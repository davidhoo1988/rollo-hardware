module comb_SA #(parameter DAT_W = 101)(
  input wire clk,
  input wire rst_b,
  input wire mode,
  input start,
  input wire [DAT_W-1:0] data,
  output reg finish,
  output wire full_rank,
  output wire [DAT_W-1:0] result
);

  reg [5 : 1] start_tmp;
  reg [5 : 1] start_row;

  always @(posedge clk) begin
    start_tmp[1] <= start;
    start_row[1] <= start_tmp[1];
    start_tmp[2] <= start_row[1];
    start_row[2] <= start_tmp[2];
    start_tmp[3] <= start_row[2];
    start_row[3] <= start_tmp[3];
    start_tmp[4] <= start_row[3];
    start_row[4] <= start_tmp[4];
    start_tmp[5] <= start_row[4];
    start_row[5] <= start_tmp[5];
  end

 //input skewed form
 wire data_col0;
 reg [1:1] data_col1;
 reg [2:1] data_col2;
 reg [3:1] data_col3;
 reg [4:1] data_col4;
 reg [5:1] data_col5;
 reg [6:1] data_col6;
 reg [7:1] data_col7;
 reg [8:1] data_col8;
 reg [9:1] data_col9;
 reg [10:1] data_col10;
 reg [11:1] data_col11;
 reg [12:1] data_col12;
 reg [13:1] data_col13;
 reg [14:1] data_col14;
 reg [15:1] data_col15;
 reg [16:1] data_col16;
 reg [17:1] data_col17;
 reg [18:1] data_col18;
 reg [19:1] data_col19;
 reg [20:1] data_col20;
 reg [21:1] data_col21;
 reg [22:1] data_col22;
 reg [23:1] data_col23;
 reg [24:1] data_col24;
 reg [25:1] data_col25;
 reg [26:1] data_col26;
 reg [27:1] data_col27;
 reg [28:1] data_col28;
 reg [29:1] data_col29;
 reg [30:1] data_col30;
 reg [31:1] data_col31;
 reg [32:1] data_col32;
 reg [33:1] data_col33;
 reg [34:1] data_col34;
 reg [35:1] data_col35;
 reg [36:1] data_col36;
 reg [37:1] data_col37;
 reg [38:1] data_col38;
 reg [39:1] data_col39;
 reg [40:1] data_col40;
 reg [41:1] data_col41;
 reg [42:1] data_col42;
 reg [43:1] data_col43;
 reg [44:1] data_col44;
 reg [45:1] data_col45;
 reg [46:1] data_col46;
 reg [47:1] data_col47;
 reg [48:1] data_col48;
 reg [49:1] data_col49;
 reg [50:1] data_col50;
 reg [51:1] data_col51;
 reg [52:1] data_col52;
 reg [53:1] data_col53;
 reg [54:1] data_col54;
 reg [55:1] data_col55;
 reg [56:1] data_col56;
 reg [57:1] data_col57;
 reg [58:1] data_col58;
 reg [59:1] data_col59;
 reg [60:1] data_col60;
 reg [61:1] data_col61;
 reg [62:1] data_col62;
 reg [63:1] data_col63;
 reg [64:1] data_col64;
 reg [65:1] data_col65;
 reg [66:1] data_col66;
 reg [67:1] data_col67;
 reg [68:1] data_col68;
 reg [69:1] data_col69;
 reg [70:1] data_col70;
 reg [71:1] data_col71;
 reg [72:1] data_col72;
 reg [73:1] data_col73;
 reg [74:1] data_col74;
 reg [75:1] data_col75;
 reg [76:1] data_col76;
 reg [77:1] data_col77;
 reg [78:1] data_col78;
 reg [79:1] data_col79;
 reg [80:1] data_col80;
 reg [81:1] data_col81;
 reg [82:1] data_col82;
 reg [83:1] data_col83;
 reg [84:1] data_col84;
 reg [85:1] data_col85;
 reg [86:1] data_col86;
 reg [87:1] data_col87;
 reg [88:1] data_col88;
 reg [89:1] data_col89;
 reg [90:1] data_col90;
 reg [91:1] data_col91;
 reg [92:1] data_col92;
 reg [93:1] data_col93;
 reg [94:1] data_col94;
 reg [95:1] data_col95;
 reg [96:1] data_col96;
 reg [97:1] data_col97;
 reg [98:1] data_col98;
 reg [99:1] data_col99;
 reg [100:1] data_col100;

 assign data_col0 = data[100];

  always @(posedge clk) begin
   data_col1[1] <= data[99];

   data_col2[1] <= data[98];
   data_col2[2] <= data_col2[1];

   data_col3[1] <= data[97];
   data_col3[2] <= data_col3[1];
   data_col3[3] <= data_col3[2];

   data_col4[1] <= data[96];
   data_col4[2] <= data_col4[1];
   data_col4[3] <= data_col4[2];
   data_col4[4] <= data_col4[3];

   data_col5[1] <= data[95];
   data_col5[2] <= data_col5[1];
   data_col5[3] <= data_col5[2];
   data_col5[4] <= data_col5[3];
   data_col5[5] <= data_col5[4];

   data_col6[1] <= data[94];
   data_col6[2] <= data_col6[1];
   data_col6[3] <= data_col6[2];
   data_col6[4] <= data_col6[3];
   data_col6[5] <= data_col6[4];
   data_col6[6] <= data_col6[5];

   data_col7[1] <= data[93];
   data_col7[2] <= data_col7[1];
   data_col7[3] <= data_col7[2];
   data_col7[4] <= data_col7[3];
   data_col7[5] <= data_col7[4];
   data_col7[6] <= data_col7[5];
   data_col7[7] <= data_col7[6];

   data_col8[1] <= data[92];
   data_col8[2] <= data_col8[1];
   data_col8[3] <= data_col8[2];
   data_col8[4] <= data_col8[3];
   data_col8[5] <= data_col8[4];
   data_col8[6] <= data_col8[5];
   data_col8[7] <= data_col8[6];
   data_col8[8] <= data_col8[7];

   data_col9[1] <= data[91];
   data_col9[2] <= data_col9[1];
   data_col9[3] <= data_col9[2];
   data_col9[4] <= data_col9[3];
   data_col9[5] <= data_col9[4];
   data_col9[6] <= data_col9[5];
   data_col9[7] <= data_col9[6];
   data_col9[8] <= data_col9[7];
   data_col9[9] <= data_col9[8];

   data_col10[1] <= data[90];
   data_col10[2] <= data_col10[1];
   data_col10[3] <= data_col10[2];
   data_col10[4] <= data_col10[3];
   data_col10[5] <= data_col10[4];
   data_col10[6] <= data_col10[5];
   data_col10[7] <= data_col10[6];
   data_col10[8] <= data_col10[7];
   data_col10[9] <= data_col10[8];
   data_col10[10] <= data_col10[9];

   data_col11[1] <= data[89];
   data_col11[2] <= data_col11[1];
   data_col11[3] <= data_col11[2];
   data_col11[4] <= data_col11[3];
   data_col11[5] <= data_col11[4];
   data_col11[6] <= data_col11[5];
   data_col11[7] <= data_col11[6];
   data_col11[8] <= data_col11[7];
   data_col11[9] <= data_col11[8];
   data_col11[10] <= data_col11[9];
   data_col11[11] <= data_col11[10];

   data_col12[1] <= data[88];
   data_col12[2] <= data_col12[1];
   data_col12[3] <= data_col12[2];
   data_col12[4] <= data_col12[3];
   data_col12[5] <= data_col12[4];
   data_col12[6] <= data_col12[5];
   data_col12[7] <= data_col12[6];
   data_col12[8] <= data_col12[7];
   data_col12[9] <= data_col12[8];
   data_col12[10] <= data_col12[9];
   data_col12[11] <= data_col12[10];
   data_col12[12] <= data_col12[11];

   data_col13[1] <= data[87];
   data_col13[2] <= data_col13[1];
   data_col13[3] <= data_col13[2];
   data_col13[4] <= data_col13[3];
   data_col13[5] <= data_col13[4];
   data_col13[6] <= data_col13[5];
   data_col13[7] <= data_col13[6];
   data_col13[8] <= data_col13[7];
   data_col13[9] <= data_col13[8];
   data_col13[10] <= data_col13[9];
   data_col13[11] <= data_col13[10];
   data_col13[12] <= data_col13[11];
   data_col13[13] <= data_col13[12];

   data_col14[1] <= data[86];
   data_col14[2] <= data_col14[1];
   data_col14[3] <= data_col14[2];
   data_col14[4] <= data_col14[3];
   data_col14[5] <= data_col14[4];
   data_col14[6] <= data_col14[5];
   data_col14[7] <= data_col14[6];
   data_col14[8] <= data_col14[7];
   data_col14[9] <= data_col14[8];
   data_col14[10] <= data_col14[9];
   data_col14[11] <= data_col14[10];
   data_col14[12] <= data_col14[11];
   data_col14[13] <= data_col14[12];
   data_col14[14] <= data_col14[13];

   data_col15[1] <= data[85];
   data_col15[2] <= data_col15[1];
   data_col15[3] <= data_col15[2];
   data_col15[4] <= data_col15[3];
   data_col15[5] <= data_col15[4];
   data_col15[6] <= data_col15[5];
   data_col15[7] <= data_col15[6];
   data_col15[8] <= data_col15[7];
   data_col15[9] <= data_col15[8];
   data_col15[10] <= data_col15[9];
   data_col15[11] <= data_col15[10];
   data_col15[12] <= data_col15[11];
   data_col15[13] <= data_col15[12];
   data_col15[14] <= data_col15[13];
   data_col15[15] <= data_col15[14];

   data_col16[1] <= data[84];
   data_col16[2] <= data_col16[1];
   data_col16[3] <= data_col16[2];
   data_col16[4] <= data_col16[3];
   data_col16[5] <= data_col16[4];
   data_col16[6] <= data_col16[5];
   data_col16[7] <= data_col16[6];
   data_col16[8] <= data_col16[7];
   data_col16[9] <= data_col16[8];
   data_col16[10] <= data_col16[9];
   data_col16[11] <= data_col16[10];
   data_col16[12] <= data_col16[11];
   data_col16[13] <= data_col16[12];
   data_col16[14] <= data_col16[13];
   data_col16[15] <= data_col16[14];
   data_col16[16] <= data_col16[15];

   data_col17[1] <= data[83];
   data_col17[2] <= data_col17[1];
   data_col17[3] <= data_col17[2];
   data_col17[4] <= data_col17[3];
   data_col17[5] <= data_col17[4];
   data_col17[6] <= data_col17[5];
   data_col17[7] <= data_col17[6];
   data_col17[8] <= data_col17[7];
   data_col17[9] <= data_col17[8];
   data_col17[10] <= data_col17[9];
   data_col17[11] <= data_col17[10];
   data_col17[12] <= data_col17[11];
   data_col17[13] <= data_col17[12];
   data_col17[14] <= data_col17[13];
   data_col17[15] <= data_col17[14];
   data_col17[16] <= data_col17[15];
   data_col17[17] <= data_col17[16];

   data_col18[1] <= data[82];
   data_col18[2] <= data_col18[1];
   data_col18[3] <= data_col18[2];
   data_col18[4] <= data_col18[3];
   data_col18[5] <= data_col18[4];
   data_col18[6] <= data_col18[5];
   data_col18[7] <= data_col18[6];
   data_col18[8] <= data_col18[7];
   data_col18[9] <= data_col18[8];
   data_col18[10] <= data_col18[9];
   data_col18[11] <= data_col18[10];
   data_col18[12] <= data_col18[11];
   data_col18[13] <= data_col18[12];
   data_col18[14] <= data_col18[13];
   data_col18[15] <= data_col18[14];
   data_col18[16] <= data_col18[15];
   data_col18[17] <= data_col18[16];
   data_col18[18] <= data_col18[17];

   data_col19[1] <= data[81];
   data_col19[2] <= data_col19[1];
   data_col19[3] <= data_col19[2];
   data_col19[4] <= data_col19[3];
   data_col19[5] <= data_col19[4];
   data_col19[6] <= data_col19[5];
   data_col19[7] <= data_col19[6];
   data_col19[8] <= data_col19[7];
   data_col19[9] <= data_col19[8];
   data_col19[10] <= data_col19[9];
   data_col19[11] <= data_col19[10];
   data_col19[12] <= data_col19[11];
   data_col19[13] <= data_col19[12];
   data_col19[14] <= data_col19[13];
   data_col19[15] <= data_col19[14];
   data_col19[16] <= data_col19[15];
   data_col19[17] <= data_col19[16];
   data_col19[18] <= data_col19[17];
   data_col19[19] <= data_col19[18];

   data_col20[1] <= data[80];
   data_col20[2] <= data_col20[1];
   data_col20[3] <= data_col20[2];
   data_col20[4] <= data_col20[3];
   data_col20[5] <= data_col20[4];
   data_col20[6] <= data_col20[5];
   data_col20[7] <= data_col20[6];
   data_col20[8] <= data_col20[7];
   data_col20[9] <= data_col20[8];
   data_col20[10] <= data_col20[9];
   data_col20[11] <= data_col20[10];
   data_col20[12] <= data_col20[11];
   data_col20[13] <= data_col20[12];
   data_col20[14] <= data_col20[13];
   data_col20[15] <= data_col20[14];
   data_col20[16] <= data_col20[15];
   data_col20[17] <= data_col20[16];
   data_col20[18] <= data_col20[17];
   data_col20[19] <= data_col20[18];
   data_col20[20] <= data_col20[19];

   data_col21[1] <= data[79];
   data_col21[2] <= data_col21[1];
   data_col21[3] <= data_col21[2];
   data_col21[4] <= data_col21[3];
   data_col21[5] <= data_col21[4];
   data_col21[6] <= data_col21[5];
   data_col21[7] <= data_col21[6];
   data_col21[8] <= data_col21[7];
   data_col21[9] <= data_col21[8];
   data_col21[10] <= data_col21[9];
   data_col21[11] <= data_col21[10];
   data_col21[12] <= data_col21[11];
   data_col21[13] <= data_col21[12];
   data_col21[14] <= data_col21[13];
   data_col21[15] <= data_col21[14];
   data_col21[16] <= data_col21[15];
   data_col21[17] <= data_col21[16];
   data_col21[18] <= data_col21[17];
   data_col21[19] <= data_col21[18];
   data_col21[20] <= data_col21[19];
   data_col21[21] <= data_col21[20];

   data_col22[1] <= data[78];
   data_col22[2] <= data_col22[1];
   data_col22[3] <= data_col22[2];
   data_col22[4] <= data_col22[3];
   data_col22[5] <= data_col22[4];
   data_col22[6] <= data_col22[5];
   data_col22[7] <= data_col22[6];
   data_col22[8] <= data_col22[7];
   data_col22[9] <= data_col22[8];
   data_col22[10] <= data_col22[9];
   data_col22[11] <= data_col22[10];
   data_col22[12] <= data_col22[11];
   data_col22[13] <= data_col22[12];
   data_col22[14] <= data_col22[13];
   data_col22[15] <= data_col22[14];
   data_col22[16] <= data_col22[15];
   data_col22[17] <= data_col22[16];
   data_col22[18] <= data_col22[17];
   data_col22[19] <= data_col22[18];
   data_col22[20] <= data_col22[19];
   data_col22[21] <= data_col22[20];
   data_col22[22] <= data_col22[21];

   data_col23[1] <= data[77];
   data_col23[2] <= data_col23[1];
   data_col23[3] <= data_col23[2];
   data_col23[4] <= data_col23[3];
   data_col23[5] <= data_col23[4];
   data_col23[6] <= data_col23[5];
   data_col23[7] <= data_col23[6];
   data_col23[8] <= data_col23[7];
   data_col23[9] <= data_col23[8];
   data_col23[10] <= data_col23[9];
   data_col23[11] <= data_col23[10];
   data_col23[12] <= data_col23[11];
   data_col23[13] <= data_col23[12];
   data_col23[14] <= data_col23[13];
   data_col23[15] <= data_col23[14];
   data_col23[16] <= data_col23[15];
   data_col23[17] <= data_col23[16];
   data_col23[18] <= data_col23[17];
   data_col23[19] <= data_col23[18];
   data_col23[20] <= data_col23[19];
   data_col23[21] <= data_col23[20];
   data_col23[22] <= data_col23[21];
   data_col23[23] <= data_col23[22];

   data_col24[1] <= data[76];
   data_col24[2] <= data_col24[1];
   data_col24[3] <= data_col24[2];
   data_col24[4] <= data_col24[3];
   data_col24[5] <= data_col24[4];
   data_col24[6] <= data_col24[5];
   data_col24[7] <= data_col24[6];
   data_col24[8] <= data_col24[7];
   data_col24[9] <= data_col24[8];
   data_col24[10] <= data_col24[9];
   data_col24[11] <= data_col24[10];
   data_col24[12] <= data_col24[11];
   data_col24[13] <= data_col24[12];
   data_col24[14] <= data_col24[13];
   data_col24[15] <= data_col24[14];
   data_col24[16] <= data_col24[15];
   data_col24[17] <= data_col24[16];
   data_col24[18] <= data_col24[17];
   data_col24[19] <= data_col24[18];
   data_col24[20] <= data_col24[19];
   data_col24[21] <= data_col24[20];
   data_col24[22] <= data_col24[21];
   data_col24[23] <= data_col24[22];
   data_col24[24] <= data_col24[23];

   data_col25[1] <= data[75];
   data_col25[2] <= data_col25[1];
   data_col25[3] <= data_col25[2];
   data_col25[4] <= data_col25[3];
   data_col25[5] <= data_col25[4];
   data_col25[6] <= data_col25[5];
   data_col25[7] <= data_col25[6];
   data_col25[8] <= data_col25[7];
   data_col25[9] <= data_col25[8];
   data_col25[10] <= data_col25[9];
   data_col25[11] <= data_col25[10];
   data_col25[12] <= data_col25[11];
   data_col25[13] <= data_col25[12];
   data_col25[14] <= data_col25[13];
   data_col25[15] <= data_col25[14];
   data_col25[16] <= data_col25[15];
   data_col25[17] <= data_col25[16];
   data_col25[18] <= data_col25[17];
   data_col25[19] <= data_col25[18];
   data_col25[20] <= data_col25[19];
   data_col25[21] <= data_col25[20];
   data_col25[22] <= data_col25[21];
   data_col25[23] <= data_col25[22];
   data_col25[24] <= data_col25[23];
   data_col25[25] <= data_col25[24];

   data_col26[1] <= data[74];
   data_col26[2] <= data_col26[1];
   data_col26[3] <= data_col26[2];
   data_col26[4] <= data_col26[3];
   data_col26[5] <= data_col26[4];
   data_col26[6] <= data_col26[5];
   data_col26[7] <= data_col26[6];
   data_col26[8] <= data_col26[7];
   data_col26[9] <= data_col26[8];
   data_col26[10] <= data_col26[9];
   data_col26[11] <= data_col26[10];
   data_col26[12] <= data_col26[11];
   data_col26[13] <= data_col26[12];
   data_col26[14] <= data_col26[13];
   data_col26[15] <= data_col26[14];
   data_col26[16] <= data_col26[15];
   data_col26[17] <= data_col26[16];
   data_col26[18] <= data_col26[17];
   data_col26[19] <= data_col26[18];
   data_col26[20] <= data_col26[19];
   data_col26[21] <= data_col26[20];
   data_col26[22] <= data_col26[21];
   data_col26[23] <= data_col26[22];
   data_col26[24] <= data_col26[23];
   data_col26[25] <= data_col26[24];
   data_col26[26] <= data_col26[25];

   data_col27[1] <= data[73];
   data_col27[2] <= data_col27[1];
   data_col27[3] <= data_col27[2];
   data_col27[4] <= data_col27[3];
   data_col27[5] <= data_col27[4];
   data_col27[6] <= data_col27[5];
   data_col27[7] <= data_col27[6];
   data_col27[8] <= data_col27[7];
   data_col27[9] <= data_col27[8];
   data_col27[10] <= data_col27[9];
   data_col27[11] <= data_col27[10];
   data_col27[12] <= data_col27[11];
   data_col27[13] <= data_col27[12];
   data_col27[14] <= data_col27[13];
   data_col27[15] <= data_col27[14];
   data_col27[16] <= data_col27[15];
   data_col27[17] <= data_col27[16];
   data_col27[18] <= data_col27[17];
   data_col27[19] <= data_col27[18];
   data_col27[20] <= data_col27[19];
   data_col27[21] <= data_col27[20];
   data_col27[22] <= data_col27[21];
   data_col27[23] <= data_col27[22];
   data_col27[24] <= data_col27[23];
   data_col27[25] <= data_col27[24];
   data_col27[26] <= data_col27[25];
   data_col27[27] <= data_col27[26];

   data_col28[1] <= data[72];
   data_col28[2] <= data_col28[1];
   data_col28[3] <= data_col28[2];
   data_col28[4] <= data_col28[3];
   data_col28[5] <= data_col28[4];
   data_col28[6] <= data_col28[5];
   data_col28[7] <= data_col28[6];
   data_col28[8] <= data_col28[7];
   data_col28[9] <= data_col28[8];
   data_col28[10] <= data_col28[9];
   data_col28[11] <= data_col28[10];
   data_col28[12] <= data_col28[11];
   data_col28[13] <= data_col28[12];
   data_col28[14] <= data_col28[13];
   data_col28[15] <= data_col28[14];
   data_col28[16] <= data_col28[15];
   data_col28[17] <= data_col28[16];
   data_col28[18] <= data_col28[17];
   data_col28[19] <= data_col28[18];
   data_col28[20] <= data_col28[19];
   data_col28[21] <= data_col28[20];
   data_col28[22] <= data_col28[21];
   data_col28[23] <= data_col28[22];
   data_col28[24] <= data_col28[23];
   data_col28[25] <= data_col28[24];
   data_col28[26] <= data_col28[25];
   data_col28[27] <= data_col28[26];
   data_col28[28] <= data_col28[27];

   data_col29[1] <= data[71];
   data_col29[2] <= data_col29[1];
   data_col29[3] <= data_col29[2];
   data_col29[4] <= data_col29[3];
   data_col29[5] <= data_col29[4];
   data_col29[6] <= data_col29[5];
   data_col29[7] <= data_col29[6];
   data_col29[8] <= data_col29[7];
   data_col29[9] <= data_col29[8];
   data_col29[10] <= data_col29[9];
   data_col29[11] <= data_col29[10];
   data_col29[12] <= data_col29[11];
   data_col29[13] <= data_col29[12];
   data_col29[14] <= data_col29[13];
   data_col29[15] <= data_col29[14];
   data_col29[16] <= data_col29[15];
   data_col29[17] <= data_col29[16];
   data_col29[18] <= data_col29[17];
   data_col29[19] <= data_col29[18];
   data_col29[20] <= data_col29[19];
   data_col29[21] <= data_col29[20];
   data_col29[22] <= data_col29[21];
   data_col29[23] <= data_col29[22];
   data_col29[24] <= data_col29[23];
   data_col29[25] <= data_col29[24];
   data_col29[26] <= data_col29[25];
   data_col29[27] <= data_col29[26];
   data_col29[28] <= data_col29[27];
   data_col29[29] <= data_col29[28];

   data_col30[1] <= data[70];
   data_col30[2] <= data_col30[1];
   data_col30[3] <= data_col30[2];
   data_col30[4] <= data_col30[3];
   data_col30[5] <= data_col30[4];
   data_col30[6] <= data_col30[5];
   data_col30[7] <= data_col30[6];
   data_col30[8] <= data_col30[7];
   data_col30[9] <= data_col30[8];
   data_col30[10] <= data_col30[9];
   data_col30[11] <= data_col30[10];
   data_col30[12] <= data_col30[11];
   data_col30[13] <= data_col30[12];
   data_col30[14] <= data_col30[13];
   data_col30[15] <= data_col30[14];
   data_col30[16] <= data_col30[15];
   data_col30[17] <= data_col30[16];
   data_col30[18] <= data_col30[17];
   data_col30[19] <= data_col30[18];
   data_col30[20] <= data_col30[19];
   data_col30[21] <= data_col30[20];
   data_col30[22] <= data_col30[21];
   data_col30[23] <= data_col30[22];
   data_col30[24] <= data_col30[23];
   data_col30[25] <= data_col30[24];
   data_col30[26] <= data_col30[25];
   data_col30[27] <= data_col30[26];
   data_col30[28] <= data_col30[27];
   data_col30[29] <= data_col30[28];
   data_col30[30] <= data_col30[29];

   data_col31[1] <= data[69];
   data_col31[2] <= data_col31[1];
   data_col31[3] <= data_col31[2];
   data_col31[4] <= data_col31[3];
   data_col31[5] <= data_col31[4];
   data_col31[6] <= data_col31[5];
   data_col31[7] <= data_col31[6];
   data_col31[8] <= data_col31[7];
   data_col31[9] <= data_col31[8];
   data_col31[10] <= data_col31[9];
   data_col31[11] <= data_col31[10];
   data_col31[12] <= data_col31[11];
   data_col31[13] <= data_col31[12];
   data_col31[14] <= data_col31[13];
   data_col31[15] <= data_col31[14];
   data_col31[16] <= data_col31[15];
   data_col31[17] <= data_col31[16];
   data_col31[18] <= data_col31[17];
   data_col31[19] <= data_col31[18];
   data_col31[20] <= data_col31[19];
   data_col31[21] <= data_col31[20];
   data_col31[22] <= data_col31[21];
   data_col31[23] <= data_col31[22];
   data_col31[24] <= data_col31[23];
   data_col31[25] <= data_col31[24];
   data_col31[26] <= data_col31[25];
   data_col31[27] <= data_col31[26];
   data_col31[28] <= data_col31[27];
   data_col31[29] <= data_col31[28];
   data_col31[30] <= data_col31[29];
   data_col31[31] <= data_col31[30];

   data_col32[1] <= data[68];
   data_col32[2] <= data_col32[1];
   data_col32[3] <= data_col32[2];
   data_col32[4] <= data_col32[3];
   data_col32[5] <= data_col32[4];
   data_col32[6] <= data_col32[5];
   data_col32[7] <= data_col32[6];
   data_col32[8] <= data_col32[7];
   data_col32[9] <= data_col32[8];
   data_col32[10] <= data_col32[9];
   data_col32[11] <= data_col32[10];
   data_col32[12] <= data_col32[11];
   data_col32[13] <= data_col32[12];
   data_col32[14] <= data_col32[13];
   data_col32[15] <= data_col32[14];
   data_col32[16] <= data_col32[15];
   data_col32[17] <= data_col32[16];
   data_col32[18] <= data_col32[17];
   data_col32[19] <= data_col32[18];
   data_col32[20] <= data_col32[19];
   data_col32[21] <= data_col32[20];
   data_col32[22] <= data_col32[21];
   data_col32[23] <= data_col32[22];
   data_col32[24] <= data_col32[23];
   data_col32[25] <= data_col32[24];
   data_col32[26] <= data_col32[25];
   data_col32[27] <= data_col32[26];
   data_col32[28] <= data_col32[27];
   data_col32[29] <= data_col32[28];
   data_col32[30] <= data_col32[29];
   data_col32[31] <= data_col32[30];
   data_col32[32] <= data_col32[31];

   data_col33[1] <= data[67];
   data_col33[2] <= data_col33[1];
   data_col33[3] <= data_col33[2];
   data_col33[4] <= data_col33[3];
   data_col33[5] <= data_col33[4];
   data_col33[6] <= data_col33[5];
   data_col33[7] <= data_col33[6];
   data_col33[8] <= data_col33[7];
   data_col33[9] <= data_col33[8];
   data_col33[10] <= data_col33[9];
   data_col33[11] <= data_col33[10];
   data_col33[12] <= data_col33[11];
   data_col33[13] <= data_col33[12];
   data_col33[14] <= data_col33[13];
   data_col33[15] <= data_col33[14];
   data_col33[16] <= data_col33[15];
   data_col33[17] <= data_col33[16];
   data_col33[18] <= data_col33[17];
   data_col33[19] <= data_col33[18];
   data_col33[20] <= data_col33[19];
   data_col33[21] <= data_col33[20];
   data_col33[22] <= data_col33[21];
   data_col33[23] <= data_col33[22];
   data_col33[24] <= data_col33[23];
   data_col33[25] <= data_col33[24];
   data_col33[26] <= data_col33[25];
   data_col33[27] <= data_col33[26];
   data_col33[28] <= data_col33[27];
   data_col33[29] <= data_col33[28];
   data_col33[30] <= data_col33[29];
   data_col33[31] <= data_col33[30];
   data_col33[32] <= data_col33[31];
   data_col33[33] <= data_col33[32];

   data_col34[1] <= data[66];
   data_col34[2] <= data_col34[1];
   data_col34[3] <= data_col34[2];
   data_col34[4] <= data_col34[3];
   data_col34[5] <= data_col34[4];
   data_col34[6] <= data_col34[5];
   data_col34[7] <= data_col34[6];
   data_col34[8] <= data_col34[7];
   data_col34[9] <= data_col34[8];
   data_col34[10] <= data_col34[9];
   data_col34[11] <= data_col34[10];
   data_col34[12] <= data_col34[11];
   data_col34[13] <= data_col34[12];
   data_col34[14] <= data_col34[13];
   data_col34[15] <= data_col34[14];
   data_col34[16] <= data_col34[15];
   data_col34[17] <= data_col34[16];
   data_col34[18] <= data_col34[17];
   data_col34[19] <= data_col34[18];
   data_col34[20] <= data_col34[19];
   data_col34[21] <= data_col34[20];
   data_col34[22] <= data_col34[21];
   data_col34[23] <= data_col34[22];
   data_col34[24] <= data_col34[23];
   data_col34[25] <= data_col34[24];
   data_col34[26] <= data_col34[25];
   data_col34[27] <= data_col34[26];
   data_col34[28] <= data_col34[27];
   data_col34[29] <= data_col34[28];
   data_col34[30] <= data_col34[29];
   data_col34[31] <= data_col34[30];
   data_col34[32] <= data_col34[31];
   data_col34[33] <= data_col34[32];
   data_col34[34] <= data_col34[33];

   data_col35[1] <= data[65];
   data_col35[2] <= data_col35[1];
   data_col35[3] <= data_col35[2];
   data_col35[4] <= data_col35[3];
   data_col35[5] <= data_col35[4];
   data_col35[6] <= data_col35[5];
   data_col35[7] <= data_col35[6];
   data_col35[8] <= data_col35[7];
   data_col35[9] <= data_col35[8];
   data_col35[10] <= data_col35[9];
   data_col35[11] <= data_col35[10];
   data_col35[12] <= data_col35[11];
   data_col35[13] <= data_col35[12];
   data_col35[14] <= data_col35[13];
   data_col35[15] <= data_col35[14];
   data_col35[16] <= data_col35[15];
   data_col35[17] <= data_col35[16];
   data_col35[18] <= data_col35[17];
   data_col35[19] <= data_col35[18];
   data_col35[20] <= data_col35[19];
   data_col35[21] <= data_col35[20];
   data_col35[22] <= data_col35[21];
   data_col35[23] <= data_col35[22];
   data_col35[24] <= data_col35[23];
   data_col35[25] <= data_col35[24];
   data_col35[26] <= data_col35[25];
   data_col35[27] <= data_col35[26];
   data_col35[28] <= data_col35[27];
   data_col35[29] <= data_col35[28];
   data_col35[30] <= data_col35[29];
   data_col35[31] <= data_col35[30];
   data_col35[32] <= data_col35[31];
   data_col35[33] <= data_col35[32];
   data_col35[34] <= data_col35[33];
   data_col35[35] <= data_col35[34];

   data_col36[1] <= data[64];
   data_col36[2] <= data_col36[1];
   data_col36[3] <= data_col36[2];
   data_col36[4] <= data_col36[3];
   data_col36[5] <= data_col36[4];
   data_col36[6] <= data_col36[5];
   data_col36[7] <= data_col36[6];
   data_col36[8] <= data_col36[7];
   data_col36[9] <= data_col36[8];
   data_col36[10] <= data_col36[9];
   data_col36[11] <= data_col36[10];
   data_col36[12] <= data_col36[11];
   data_col36[13] <= data_col36[12];
   data_col36[14] <= data_col36[13];
   data_col36[15] <= data_col36[14];
   data_col36[16] <= data_col36[15];
   data_col36[17] <= data_col36[16];
   data_col36[18] <= data_col36[17];
   data_col36[19] <= data_col36[18];
   data_col36[20] <= data_col36[19];
   data_col36[21] <= data_col36[20];
   data_col36[22] <= data_col36[21];
   data_col36[23] <= data_col36[22];
   data_col36[24] <= data_col36[23];
   data_col36[25] <= data_col36[24];
   data_col36[26] <= data_col36[25];
   data_col36[27] <= data_col36[26];
   data_col36[28] <= data_col36[27];
   data_col36[29] <= data_col36[28];
   data_col36[30] <= data_col36[29];
   data_col36[31] <= data_col36[30];
   data_col36[32] <= data_col36[31];
   data_col36[33] <= data_col36[32];
   data_col36[34] <= data_col36[33];
   data_col36[35] <= data_col36[34];
   data_col36[36] <= data_col36[35];

   data_col37[1] <= data[63];
   data_col37[2] <= data_col37[1];
   data_col37[3] <= data_col37[2];
   data_col37[4] <= data_col37[3];
   data_col37[5] <= data_col37[4];
   data_col37[6] <= data_col37[5];
   data_col37[7] <= data_col37[6];
   data_col37[8] <= data_col37[7];
   data_col37[9] <= data_col37[8];
   data_col37[10] <= data_col37[9];
   data_col37[11] <= data_col37[10];
   data_col37[12] <= data_col37[11];
   data_col37[13] <= data_col37[12];
   data_col37[14] <= data_col37[13];
   data_col37[15] <= data_col37[14];
   data_col37[16] <= data_col37[15];
   data_col37[17] <= data_col37[16];
   data_col37[18] <= data_col37[17];
   data_col37[19] <= data_col37[18];
   data_col37[20] <= data_col37[19];
   data_col37[21] <= data_col37[20];
   data_col37[22] <= data_col37[21];
   data_col37[23] <= data_col37[22];
   data_col37[24] <= data_col37[23];
   data_col37[25] <= data_col37[24];
   data_col37[26] <= data_col37[25];
   data_col37[27] <= data_col37[26];
   data_col37[28] <= data_col37[27];
   data_col37[29] <= data_col37[28];
   data_col37[30] <= data_col37[29];
   data_col37[31] <= data_col37[30];
   data_col37[32] <= data_col37[31];
   data_col37[33] <= data_col37[32];
   data_col37[34] <= data_col37[33];
   data_col37[35] <= data_col37[34];
   data_col37[36] <= data_col37[35];
   data_col37[37] <= data_col37[36];

   data_col38[1] <= data[62];
   data_col38[2] <= data_col38[1];
   data_col38[3] <= data_col38[2];
   data_col38[4] <= data_col38[3];
   data_col38[5] <= data_col38[4];
   data_col38[6] <= data_col38[5];
   data_col38[7] <= data_col38[6];
   data_col38[8] <= data_col38[7];
   data_col38[9] <= data_col38[8];
   data_col38[10] <= data_col38[9];
   data_col38[11] <= data_col38[10];
   data_col38[12] <= data_col38[11];
   data_col38[13] <= data_col38[12];
   data_col38[14] <= data_col38[13];
   data_col38[15] <= data_col38[14];
   data_col38[16] <= data_col38[15];
   data_col38[17] <= data_col38[16];
   data_col38[18] <= data_col38[17];
   data_col38[19] <= data_col38[18];
   data_col38[20] <= data_col38[19];
   data_col38[21] <= data_col38[20];
   data_col38[22] <= data_col38[21];
   data_col38[23] <= data_col38[22];
   data_col38[24] <= data_col38[23];
   data_col38[25] <= data_col38[24];
   data_col38[26] <= data_col38[25];
   data_col38[27] <= data_col38[26];
   data_col38[28] <= data_col38[27];
   data_col38[29] <= data_col38[28];
   data_col38[30] <= data_col38[29];
   data_col38[31] <= data_col38[30];
   data_col38[32] <= data_col38[31];
   data_col38[33] <= data_col38[32];
   data_col38[34] <= data_col38[33];
   data_col38[35] <= data_col38[34];
   data_col38[36] <= data_col38[35];
   data_col38[37] <= data_col38[36];
   data_col38[38] <= data_col38[37];

   data_col39[1] <= data[61];
   data_col39[2] <= data_col39[1];
   data_col39[3] <= data_col39[2];
   data_col39[4] <= data_col39[3];
   data_col39[5] <= data_col39[4];
   data_col39[6] <= data_col39[5];
   data_col39[7] <= data_col39[6];
   data_col39[8] <= data_col39[7];
   data_col39[9] <= data_col39[8];
   data_col39[10] <= data_col39[9];
   data_col39[11] <= data_col39[10];
   data_col39[12] <= data_col39[11];
   data_col39[13] <= data_col39[12];
   data_col39[14] <= data_col39[13];
   data_col39[15] <= data_col39[14];
   data_col39[16] <= data_col39[15];
   data_col39[17] <= data_col39[16];
   data_col39[18] <= data_col39[17];
   data_col39[19] <= data_col39[18];
   data_col39[20] <= data_col39[19];
   data_col39[21] <= data_col39[20];
   data_col39[22] <= data_col39[21];
   data_col39[23] <= data_col39[22];
   data_col39[24] <= data_col39[23];
   data_col39[25] <= data_col39[24];
   data_col39[26] <= data_col39[25];
   data_col39[27] <= data_col39[26];
   data_col39[28] <= data_col39[27];
   data_col39[29] <= data_col39[28];
   data_col39[30] <= data_col39[29];
   data_col39[31] <= data_col39[30];
   data_col39[32] <= data_col39[31];
   data_col39[33] <= data_col39[32];
   data_col39[34] <= data_col39[33];
   data_col39[35] <= data_col39[34];
   data_col39[36] <= data_col39[35];
   data_col39[37] <= data_col39[36];
   data_col39[38] <= data_col39[37];
   data_col39[39] <= data_col39[38];

   data_col40[1] <= data[60];
   data_col40[2] <= data_col40[1];
   data_col40[3] <= data_col40[2];
   data_col40[4] <= data_col40[3];
   data_col40[5] <= data_col40[4];
   data_col40[6] <= data_col40[5];
   data_col40[7] <= data_col40[6];
   data_col40[8] <= data_col40[7];
   data_col40[9] <= data_col40[8];
   data_col40[10] <= data_col40[9];
   data_col40[11] <= data_col40[10];
   data_col40[12] <= data_col40[11];
   data_col40[13] <= data_col40[12];
   data_col40[14] <= data_col40[13];
   data_col40[15] <= data_col40[14];
   data_col40[16] <= data_col40[15];
   data_col40[17] <= data_col40[16];
   data_col40[18] <= data_col40[17];
   data_col40[19] <= data_col40[18];
   data_col40[20] <= data_col40[19];
   data_col40[21] <= data_col40[20];
   data_col40[22] <= data_col40[21];
   data_col40[23] <= data_col40[22];
   data_col40[24] <= data_col40[23];
   data_col40[25] <= data_col40[24];
   data_col40[26] <= data_col40[25];
   data_col40[27] <= data_col40[26];
   data_col40[28] <= data_col40[27];
   data_col40[29] <= data_col40[28];
   data_col40[30] <= data_col40[29];
   data_col40[31] <= data_col40[30];
   data_col40[32] <= data_col40[31];
   data_col40[33] <= data_col40[32];
   data_col40[34] <= data_col40[33];
   data_col40[35] <= data_col40[34];
   data_col40[36] <= data_col40[35];
   data_col40[37] <= data_col40[36];
   data_col40[38] <= data_col40[37];
   data_col40[39] <= data_col40[38];
   data_col40[40] <= data_col40[39];

   data_col41[1] <= data[59];
   data_col41[2] <= data_col41[1];
   data_col41[3] <= data_col41[2];
   data_col41[4] <= data_col41[3];
   data_col41[5] <= data_col41[4];
   data_col41[6] <= data_col41[5];
   data_col41[7] <= data_col41[6];
   data_col41[8] <= data_col41[7];
   data_col41[9] <= data_col41[8];
   data_col41[10] <= data_col41[9];
   data_col41[11] <= data_col41[10];
   data_col41[12] <= data_col41[11];
   data_col41[13] <= data_col41[12];
   data_col41[14] <= data_col41[13];
   data_col41[15] <= data_col41[14];
   data_col41[16] <= data_col41[15];
   data_col41[17] <= data_col41[16];
   data_col41[18] <= data_col41[17];
   data_col41[19] <= data_col41[18];
   data_col41[20] <= data_col41[19];
   data_col41[21] <= data_col41[20];
   data_col41[22] <= data_col41[21];
   data_col41[23] <= data_col41[22];
   data_col41[24] <= data_col41[23];
   data_col41[25] <= data_col41[24];
   data_col41[26] <= data_col41[25];
   data_col41[27] <= data_col41[26];
   data_col41[28] <= data_col41[27];
   data_col41[29] <= data_col41[28];
   data_col41[30] <= data_col41[29];
   data_col41[31] <= data_col41[30];
   data_col41[32] <= data_col41[31];
   data_col41[33] <= data_col41[32];
   data_col41[34] <= data_col41[33];
   data_col41[35] <= data_col41[34];
   data_col41[36] <= data_col41[35];
   data_col41[37] <= data_col41[36];
   data_col41[38] <= data_col41[37];
   data_col41[39] <= data_col41[38];
   data_col41[40] <= data_col41[39];
   data_col41[41] <= data_col41[40];

   data_col42[1] <= data[58];
   data_col42[2] <= data_col42[1];
   data_col42[3] <= data_col42[2];
   data_col42[4] <= data_col42[3];
   data_col42[5] <= data_col42[4];
   data_col42[6] <= data_col42[5];
   data_col42[7] <= data_col42[6];
   data_col42[8] <= data_col42[7];
   data_col42[9] <= data_col42[8];
   data_col42[10] <= data_col42[9];
   data_col42[11] <= data_col42[10];
   data_col42[12] <= data_col42[11];
   data_col42[13] <= data_col42[12];
   data_col42[14] <= data_col42[13];
   data_col42[15] <= data_col42[14];
   data_col42[16] <= data_col42[15];
   data_col42[17] <= data_col42[16];
   data_col42[18] <= data_col42[17];
   data_col42[19] <= data_col42[18];
   data_col42[20] <= data_col42[19];
   data_col42[21] <= data_col42[20];
   data_col42[22] <= data_col42[21];
   data_col42[23] <= data_col42[22];
   data_col42[24] <= data_col42[23];
   data_col42[25] <= data_col42[24];
   data_col42[26] <= data_col42[25];
   data_col42[27] <= data_col42[26];
   data_col42[28] <= data_col42[27];
   data_col42[29] <= data_col42[28];
   data_col42[30] <= data_col42[29];
   data_col42[31] <= data_col42[30];
   data_col42[32] <= data_col42[31];
   data_col42[33] <= data_col42[32];
   data_col42[34] <= data_col42[33];
   data_col42[35] <= data_col42[34];
   data_col42[36] <= data_col42[35];
   data_col42[37] <= data_col42[36];
   data_col42[38] <= data_col42[37];
   data_col42[39] <= data_col42[38];
   data_col42[40] <= data_col42[39];
   data_col42[41] <= data_col42[40];
   data_col42[42] <= data_col42[41];

   data_col43[1] <= data[57];
   data_col43[2] <= data_col43[1];
   data_col43[3] <= data_col43[2];
   data_col43[4] <= data_col43[3];
   data_col43[5] <= data_col43[4];
   data_col43[6] <= data_col43[5];
   data_col43[7] <= data_col43[6];
   data_col43[8] <= data_col43[7];
   data_col43[9] <= data_col43[8];
   data_col43[10] <= data_col43[9];
   data_col43[11] <= data_col43[10];
   data_col43[12] <= data_col43[11];
   data_col43[13] <= data_col43[12];
   data_col43[14] <= data_col43[13];
   data_col43[15] <= data_col43[14];
   data_col43[16] <= data_col43[15];
   data_col43[17] <= data_col43[16];
   data_col43[18] <= data_col43[17];
   data_col43[19] <= data_col43[18];
   data_col43[20] <= data_col43[19];
   data_col43[21] <= data_col43[20];
   data_col43[22] <= data_col43[21];
   data_col43[23] <= data_col43[22];
   data_col43[24] <= data_col43[23];
   data_col43[25] <= data_col43[24];
   data_col43[26] <= data_col43[25];
   data_col43[27] <= data_col43[26];
   data_col43[28] <= data_col43[27];
   data_col43[29] <= data_col43[28];
   data_col43[30] <= data_col43[29];
   data_col43[31] <= data_col43[30];
   data_col43[32] <= data_col43[31];
   data_col43[33] <= data_col43[32];
   data_col43[34] <= data_col43[33];
   data_col43[35] <= data_col43[34];
   data_col43[36] <= data_col43[35];
   data_col43[37] <= data_col43[36];
   data_col43[38] <= data_col43[37];
   data_col43[39] <= data_col43[38];
   data_col43[40] <= data_col43[39];
   data_col43[41] <= data_col43[40];
   data_col43[42] <= data_col43[41];
   data_col43[43] <= data_col43[42];

   data_col44[1] <= data[56];
   data_col44[2] <= data_col44[1];
   data_col44[3] <= data_col44[2];
   data_col44[4] <= data_col44[3];
   data_col44[5] <= data_col44[4];
   data_col44[6] <= data_col44[5];
   data_col44[7] <= data_col44[6];
   data_col44[8] <= data_col44[7];
   data_col44[9] <= data_col44[8];
   data_col44[10] <= data_col44[9];
   data_col44[11] <= data_col44[10];
   data_col44[12] <= data_col44[11];
   data_col44[13] <= data_col44[12];
   data_col44[14] <= data_col44[13];
   data_col44[15] <= data_col44[14];
   data_col44[16] <= data_col44[15];
   data_col44[17] <= data_col44[16];
   data_col44[18] <= data_col44[17];
   data_col44[19] <= data_col44[18];
   data_col44[20] <= data_col44[19];
   data_col44[21] <= data_col44[20];
   data_col44[22] <= data_col44[21];
   data_col44[23] <= data_col44[22];
   data_col44[24] <= data_col44[23];
   data_col44[25] <= data_col44[24];
   data_col44[26] <= data_col44[25];
   data_col44[27] <= data_col44[26];
   data_col44[28] <= data_col44[27];
   data_col44[29] <= data_col44[28];
   data_col44[30] <= data_col44[29];
   data_col44[31] <= data_col44[30];
   data_col44[32] <= data_col44[31];
   data_col44[33] <= data_col44[32];
   data_col44[34] <= data_col44[33];
   data_col44[35] <= data_col44[34];
   data_col44[36] <= data_col44[35];
   data_col44[37] <= data_col44[36];
   data_col44[38] <= data_col44[37];
   data_col44[39] <= data_col44[38];
   data_col44[40] <= data_col44[39];
   data_col44[41] <= data_col44[40];
   data_col44[42] <= data_col44[41];
   data_col44[43] <= data_col44[42];
   data_col44[44] <= data_col44[43];

   data_col45[1] <= data[55];
   data_col45[2] <= data_col45[1];
   data_col45[3] <= data_col45[2];
   data_col45[4] <= data_col45[3];
   data_col45[5] <= data_col45[4];
   data_col45[6] <= data_col45[5];
   data_col45[7] <= data_col45[6];
   data_col45[8] <= data_col45[7];
   data_col45[9] <= data_col45[8];
   data_col45[10] <= data_col45[9];
   data_col45[11] <= data_col45[10];
   data_col45[12] <= data_col45[11];
   data_col45[13] <= data_col45[12];
   data_col45[14] <= data_col45[13];
   data_col45[15] <= data_col45[14];
   data_col45[16] <= data_col45[15];
   data_col45[17] <= data_col45[16];
   data_col45[18] <= data_col45[17];
   data_col45[19] <= data_col45[18];
   data_col45[20] <= data_col45[19];
   data_col45[21] <= data_col45[20];
   data_col45[22] <= data_col45[21];
   data_col45[23] <= data_col45[22];
   data_col45[24] <= data_col45[23];
   data_col45[25] <= data_col45[24];
   data_col45[26] <= data_col45[25];
   data_col45[27] <= data_col45[26];
   data_col45[28] <= data_col45[27];
   data_col45[29] <= data_col45[28];
   data_col45[30] <= data_col45[29];
   data_col45[31] <= data_col45[30];
   data_col45[32] <= data_col45[31];
   data_col45[33] <= data_col45[32];
   data_col45[34] <= data_col45[33];
   data_col45[35] <= data_col45[34];
   data_col45[36] <= data_col45[35];
   data_col45[37] <= data_col45[36];
   data_col45[38] <= data_col45[37];
   data_col45[39] <= data_col45[38];
   data_col45[40] <= data_col45[39];
   data_col45[41] <= data_col45[40];
   data_col45[42] <= data_col45[41];
   data_col45[43] <= data_col45[42];
   data_col45[44] <= data_col45[43];
   data_col45[45] <= data_col45[44];

   data_col46[1] <= data[54];
   data_col46[2] <= data_col46[1];
   data_col46[3] <= data_col46[2];
   data_col46[4] <= data_col46[3];
   data_col46[5] <= data_col46[4];
   data_col46[6] <= data_col46[5];
   data_col46[7] <= data_col46[6];
   data_col46[8] <= data_col46[7];
   data_col46[9] <= data_col46[8];
   data_col46[10] <= data_col46[9];
   data_col46[11] <= data_col46[10];
   data_col46[12] <= data_col46[11];
   data_col46[13] <= data_col46[12];
   data_col46[14] <= data_col46[13];
   data_col46[15] <= data_col46[14];
   data_col46[16] <= data_col46[15];
   data_col46[17] <= data_col46[16];
   data_col46[18] <= data_col46[17];
   data_col46[19] <= data_col46[18];
   data_col46[20] <= data_col46[19];
   data_col46[21] <= data_col46[20];
   data_col46[22] <= data_col46[21];
   data_col46[23] <= data_col46[22];
   data_col46[24] <= data_col46[23];
   data_col46[25] <= data_col46[24];
   data_col46[26] <= data_col46[25];
   data_col46[27] <= data_col46[26];
   data_col46[28] <= data_col46[27];
   data_col46[29] <= data_col46[28];
   data_col46[30] <= data_col46[29];
   data_col46[31] <= data_col46[30];
   data_col46[32] <= data_col46[31];
   data_col46[33] <= data_col46[32];
   data_col46[34] <= data_col46[33];
   data_col46[35] <= data_col46[34];
   data_col46[36] <= data_col46[35];
   data_col46[37] <= data_col46[36];
   data_col46[38] <= data_col46[37];
   data_col46[39] <= data_col46[38];
   data_col46[40] <= data_col46[39];
   data_col46[41] <= data_col46[40];
   data_col46[42] <= data_col46[41];
   data_col46[43] <= data_col46[42];
   data_col46[44] <= data_col46[43];
   data_col46[45] <= data_col46[44];
   data_col46[46] <= data_col46[45];

   data_col47[1] <= data[53];
   data_col47[2] <= data_col47[1];
   data_col47[3] <= data_col47[2];
   data_col47[4] <= data_col47[3];
   data_col47[5] <= data_col47[4];
   data_col47[6] <= data_col47[5];
   data_col47[7] <= data_col47[6];
   data_col47[8] <= data_col47[7];
   data_col47[9] <= data_col47[8];
   data_col47[10] <= data_col47[9];
   data_col47[11] <= data_col47[10];
   data_col47[12] <= data_col47[11];
   data_col47[13] <= data_col47[12];
   data_col47[14] <= data_col47[13];
   data_col47[15] <= data_col47[14];
   data_col47[16] <= data_col47[15];
   data_col47[17] <= data_col47[16];
   data_col47[18] <= data_col47[17];
   data_col47[19] <= data_col47[18];
   data_col47[20] <= data_col47[19];
   data_col47[21] <= data_col47[20];
   data_col47[22] <= data_col47[21];
   data_col47[23] <= data_col47[22];
   data_col47[24] <= data_col47[23];
   data_col47[25] <= data_col47[24];
   data_col47[26] <= data_col47[25];
   data_col47[27] <= data_col47[26];
   data_col47[28] <= data_col47[27];
   data_col47[29] <= data_col47[28];
   data_col47[30] <= data_col47[29];
   data_col47[31] <= data_col47[30];
   data_col47[32] <= data_col47[31];
   data_col47[33] <= data_col47[32];
   data_col47[34] <= data_col47[33];
   data_col47[35] <= data_col47[34];
   data_col47[36] <= data_col47[35];
   data_col47[37] <= data_col47[36];
   data_col47[38] <= data_col47[37];
   data_col47[39] <= data_col47[38];
   data_col47[40] <= data_col47[39];
   data_col47[41] <= data_col47[40];
   data_col47[42] <= data_col47[41];
   data_col47[43] <= data_col47[42];
   data_col47[44] <= data_col47[43];
   data_col47[45] <= data_col47[44];
   data_col47[46] <= data_col47[45];
   data_col47[47] <= data_col47[46];

   data_col48[1] <= data[52];
   data_col48[2] <= data_col48[1];
   data_col48[3] <= data_col48[2];
   data_col48[4] <= data_col48[3];
   data_col48[5] <= data_col48[4];
   data_col48[6] <= data_col48[5];
   data_col48[7] <= data_col48[6];
   data_col48[8] <= data_col48[7];
   data_col48[9] <= data_col48[8];
   data_col48[10] <= data_col48[9];
   data_col48[11] <= data_col48[10];
   data_col48[12] <= data_col48[11];
   data_col48[13] <= data_col48[12];
   data_col48[14] <= data_col48[13];
   data_col48[15] <= data_col48[14];
   data_col48[16] <= data_col48[15];
   data_col48[17] <= data_col48[16];
   data_col48[18] <= data_col48[17];
   data_col48[19] <= data_col48[18];
   data_col48[20] <= data_col48[19];
   data_col48[21] <= data_col48[20];
   data_col48[22] <= data_col48[21];
   data_col48[23] <= data_col48[22];
   data_col48[24] <= data_col48[23];
   data_col48[25] <= data_col48[24];
   data_col48[26] <= data_col48[25];
   data_col48[27] <= data_col48[26];
   data_col48[28] <= data_col48[27];
   data_col48[29] <= data_col48[28];
   data_col48[30] <= data_col48[29];
   data_col48[31] <= data_col48[30];
   data_col48[32] <= data_col48[31];
   data_col48[33] <= data_col48[32];
   data_col48[34] <= data_col48[33];
   data_col48[35] <= data_col48[34];
   data_col48[36] <= data_col48[35];
   data_col48[37] <= data_col48[36];
   data_col48[38] <= data_col48[37];
   data_col48[39] <= data_col48[38];
   data_col48[40] <= data_col48[39];
   data_col48[41] <= data_col48[40];
   data_col48[42] <= data_col48[41];
   data_col48[43] <= data_col48[42];
   data_col48[44] <= data_col48[43];
   data_col48[45] <= data_col48[44];
   data_col48[46] <= data_col48[45];
   data_col48[47] <= data_col48[46];
   data_col48[48] <= data_col48[47];

   data_col49[1] <= data[51];
   data_col49[2] <= data_col49[1];
   data_col49[3] <= data_col49[2];
   data_col49[4] <= data_col49[3];
   data_col49[5] <= data_col49[4];
   data_col49[6] <= data_col49[5];
   data_col49[7] <= data_col49[6];
   data_col49[8] <= data_col49[7];
   data_col49[9] <= data_col49[8];
   data_col49[10] <= data_col49[9];
   data_col49[11] <= data_col49[10];
   data_col49[12] <= data_col49[11];
   data_col49[13] <= data_col49[12];
   data_col49[14] <= data_col49[13];
   data_col49[15] <= data_col49[14];
   data_col49[16] <= data_col49[15];
   data_col49[17] <= data_col49[16];
   data_col49[18] <= data_col49[17];
   data_col49[19] <= data_col49[18];
   data_col49[20] <= data_col49[19];
   data_col49[21] <= data_col49[20];
   data_col49[22] <= data_col49[21];
   data_col49[23] <= data_col49[22];
   data_col49[24] <= data_col49[23];
   data_col49[25] <= data_col49[24];
   data_col49[26] <= data_col49[25];
   data_col49[27] <= data_col49[26];
   data_col49[28] <= data_col49[27];
   data_col49[29] <= data_col49[28];
   data_col49[30] <= data_col49[29];
   data_col49[31] <= data_col49[30];
   data_col49[32] <= data_col49[31];
   data_col49[33] <= data_col49[32];
   data_col49[34] <= data_col49[33];
   data_col49[35] <= data_col49[34];
   data_col49[36] <= data_col49[35];
   data_col49[37] <= data_col49[36];
   data_col49[38] <= data_col49[37];
   data_col49[39] <= data_col49[38];
   data_col49[40] <= data_col49[39];
   data_col49[41] <= data_col49[40];
   data_col49[42] <= data_col49[41];
   data_col49[43] <= data_col49[42];
   data_col49[44] <= data_col49[43];
   data_col49[45] <= data_col49[44];
   data_col49[46] <= data_col49[45];
   data_col49[47] <= data_col49[46];
   data_col49[48] <= data_col49[47];
   data_col49[49] <= data_col49[48];

   data_col50[1] <= data[50];
   data_col50[2] <= data_col50[1];
   data_col50[3] <= data_col50[2];
   data_col50[4] <= data_col50[3];
   data_col50[5] <= data_col50[4];
   data_col50[6] <= data_col50[5];
   data_col50[7] <= data_col50[6];
   data_col50[8] <= data_col50[7];
   data_col50[9] <= data_col50[8];
   data_col50[10] <= data_col50[9];
   data_col50[11] <= data_col50[10];
   data_col50[12] <= data_col50[11];
   data_col50[13] <= data_col50[12];
   data_col50[14] <= data_col50[13];
   data_col50[15] <= data_col50[14];
   data_col50[16] <= data_col50[15];
   data_col50[17] <= data_col50[16];
   data_col50[18] <= data_col50[17];
   data_col50[19] <= data_col50[18];
   data_col50[20] <= data_col50[19];
   data_col50[21] <= data_col50[20];
   data_col50[22] <= data_col50[21];
   data_col50[23] <= data_col50[22];
   data_col50[24] <= data_col50[23];
   data_col50[25] <= data_col50[24];
   data_col50[26] <= data_col50[25];
   data_col50[27] <= data_col50[26];
   data_col50[28] <= data_col50[27];
   data_col50[29] <= data_col50[28];
   data_col50[30] <= data_col50[29];
   data_col50[31] <= data_col50[30];
   data_col50[32] <= data_col50[31];
   data_col50[33] <= data_col50[32];
   data_col50[34] <= data_col50[33];
   data_col50[35] <= data_col50[34];
   data_col50[36] <= data_col50[35];
   data_col50[37] <= data_col50[36];
   data_col50[38] <= data_col50[37];
   data_col50[39] <= data_col50[38];
   data_col50[40] <= data_col50[39];
   data_col50[41] <= data_col50[40];
   data_col50[42] <= data_col50[41];
   data_col50[43] <= data_col50[42];
   data_col50[44] <= data_col50[43];
   data_col50[45] <= data_col50[44];
   data_col50[46] <= data_col50[45];
   data_col50[47] <= data_col50[46];
   data_col50[48] <= data_col50[47];
   data_col50[49] <= data_col50[48];
   data_col50[50] <= data_col50[49];

   data_col51[1] <= data[49];
   data_col51[2] <= data_col51[1];
   data_col51[3] <= data_col51[2];
   data_col51[4] <= data_col51[3];
   data_col51[5] <= data_col51[4];
   data_col51[6] <= data_col51[5];
   data_col51[7] <= data_col51[6];
   data_col51[8] <= data_col51[7];
   data_col51[9] <= data_col51[8];
   data_col51[10] <= data_col51[9];
   data_col51[11] <= data_col51[10];
   data_col51[12] <= data_col51[11];
   data_col51[13] <= data_col51[12];
   data_col51[14] <= data_col51[13];
   data_col51[15] <= data_col51[14];
   data_col51[16] <= data_col51[15];
   data_col51[17] <= data_col51[16];
   data_col51[18] <= data_col51[17];
   data_col51[19] <= data_col51[18];
   data_col51[20] <= data_col51[19];
   data_col51[21] <= data_col51[20];
   data_col51[22] <= data_col51[21];
   data_col51[23] <= data_col51[22];
   data_col51[24] <= data_col51[23];
   data_col51[25] <= data_col51[24];
   data_col51[26] <= data_col51[25];
   data_col51[27] <= data_col51[26];
   data_col51[28] <= data_col51[27];
   data_col51[29] <= data_col51[28];
   data_col51[30] <= data_col51[29];
   data_col51[31] <= data_col51[30];
   data_col51[32] <= data_col51[31];
   data_col51[33] <= data_col51[32];
   data_col51[34] <= data_col51[33];
   data_col51[35] <= data_col51[34];
   data_col51[36] <= data_col51[35];
   data_col51[37] <= data_col51[36];
   data_col51[38] <= data_col51[37];
   data_col51[39] <= data_col51[38];
   data_col51[40] <= data_col51[39];
   data_col51[41] <= data_col51[40];
   data_col51[42] <= data_col51[41];
   data_col51[43] <= data_col51[42];
   data_col51[44] <= data_col51[43];
   data_col51[45] <= data_col51[44];
   data_col51[46] <= data_col51[45];
   data_col51[47] <= data_col51[46];
   data_col51[48] <= data_col51[47];
   data_col51[49] <= data_col51[48];
   data_col51[50] <= data_col51[49];
   data_col51[51] <= data_col51[50];

   data_col52[1] <= data[48];
   data_col52[2] <= data_col52[1];
   data_col52[3] <= data_col52[2];
   data_col52[4] <= data_col52[3];
   data_col52[5] <= data_col52[4];
   data_col52[6] <= data_col52[5];
   data_col52[7] <= data_col52[6];
   data_col52[8] <= data_col52[7];
   data_col52[9] <= data_col52[8];
   data_col52[10] <= data_col52[9];
   data_col52[11] <= data_col52[10];
   data_col52[12] <= data_col52[11];
   data_col52[13] <= data_col52[12];
   data_col52[14] <= data_col52[13];
   data_col52[15] <= data_col52[14];
   data_col52[16] <= data_col52[15];
   data_col52[17] <= data_col52[16];
   data_col52[18] <= data_col52[17];
   data_col52[19] <= data_col52[18];
   data_col52[20] <= data_col52[19];
   data_col52[21] <= data_col52[20];
   data_col52[22] <= data_col52[21];
   data_col52[23] <= data_col52[22];
   data_col52[24] <= data_col52[23];
   data_col52[25] <= data_col52[24];
   data_col52[26] <= data_col52[25];
   data_col52[27] <= data_col52[26];
   data_col52[28] <= data_col52[27];
   data_col52[29] <= data_col52[28];
   data_col52[30] <= data_col52[29];
   data_col52[31] <= data_col52[30];
   data_col52[32] <= data_col52[31];
   data_col52[33] <= data_col52[32];
   data_col52[34] <= data_col52[33];
   data_col52[35] <= data_col52[34];
   data_col52[36] <= data_col52[35];
   data_col52[37] <= data_col52[36];
   data_col52[38] <= data_col52[37];
   data_col52[39] <= data_col52[38];
   data_col52[40] <= data_col52[39];
   data_col52[41] <= data_col52[40];
   data_col52[42] <= data_col52[41];
   data_col52[43] <= data_col52[42];
   data_col52[44] <= data_col52[43];
   data_col52[45] <= data_col52[44];
   data_col52[46] <= data_col52[45];
   data_col52[47] <= data_col52[46];
   data_col52[48] <= data_col52[47];
   data_col52[49] <= data_col52[48];
   data_col52[50] <= data_col52[49];
   data_col52[51] <= data_col52[50];
   data_col52[52] <= data_col52[51];

   data_col53[1] <= data[47];
   data_col53[2] <= data_col53[1];
   data_col53[3] <= data_col53[2];
   data_col53[4] <= data_col53[3];
   data_col53[5] <= data_col53[4];
   data_col53[6] <= data_col53[5];
   data_col53[7] <= data_col53[6];
   data_col53[8] <= data_col53[7];
   data_col53[9] <= data_col53[8];
   data_col53[10] <= data_col53[9];
   data_col53[11] <= data_col53[10];
   data_col53[12] <= data_col53[11];
   data_col53[13] <= data_col53[12];
   data_col53[14] <= data_col53[13];
   data_col53[15] <= data_col53[14];
   data_col53[16] <= data_col53[15];
   data_col53[17] <= data_col53[16];
   data_col53[18] <= data_col53[17];
   data_col53[19] <= data_col53[18];
   data_col53[20] <= data_col53[19];
   data_col53[21] <= data_col53[20];
   data_col53[22] <= data_col53[21];
   data_col53[23] <= data_col53[22];
   data_col53[24] <= data_col53[23];
   data_col53[25] <= data_col53[24];
   data_col53[26] <= data_col53[25];
   data_col53[27] <= data_col53[26];
   data_col53[28] <= data_col53[27];
   data_col53[29] <= data_col53[28];
   data_col53[30] <= data_col53[29];
   data_col53[31] <= data_col53[30];
   data_col53[32] <= data_col53[31];
   data_col53[33] <= data_col53[32];
   data_col53[34] <= data_col53[33];
   data_col53[35] <= data_col53[34];
   data_col53[36] <= data_col53[35];
   data_col53[37] <= data_col53[36];
   data_col53[38] <= data_col53[37];
   data_col53[39] <= data_col53[38];
   data_col53[40] <= data_col53[39];
   data_col53[41] <= data_col53[40];
   data_col53[42] <= data_col53[41];
   data_col53[43] <= data_col53[42];
   data_col53[44] <= data_col53[43];
   data_col53[45] <= data_col53[44];
   data_col53[46] <= data_col53[45];
   data_col53[47] <= data_col53[46];
   data_col53[48] <= data_col53[47];
   data_col53[49] <= data_col53[48];
   data_col53[50] <= data_col53[49];
   data_col53[51] <= data_col53[50];
   data_col53[52] <= data_col53[51];
   data_col53[53] <= data_col53[52];

   data_col54[1] <= data[46];
   data_col54[2] <= data_col54[1];
   data_col54[3] <= data_col54[2];
   data_col54[4] <= data_col54[3];
   data_col54[5] <= data_col54[4];
   data_col54[6] <= data_col54[5];
   data_col54[7] <= data_col54[6];
   data_col54[8] <= data_col54[7];
   data_col54[9] <= data_col54[8];
   data_col54[10] <= data_col54[9];
   data_col54[11] <= data_col54[10];
   data_col54[12] <= data_col54[11];
   data_col54[13] <= data_col54[12];
   data_col54[14] <= data_col54[13];
   data_col54[15] <= data_col54[14];
   data_col54[16] <= data_col54[15];
   data_col54[17] <= data_col54[16];
   data_col54[18] <= data_col54[17];
   data_col54[19] <= data_col54[18];
   data_col54[20] <= data_col54[19];
   data_col54[21] <= data_col54[20];
   data_col54[22] <= data_col54[21];
   data_col54[23] <= data_col54[22];
   data_col54[24] <= data_col54[23];
   data_col54[25] <= data_col54[24];
   data_col54[26] <= data_col54[25];
   data_col54[27] <= data_col54[26];
   data_col54[28] <= data_col54[27];
   data_col54[29] <= data_col54[28];
   data_col54[30] <= data_col54[29];
   data_col54[31] <= data_col54[30];
   data_col54[32] <= data_col54[31];
   data_col54[33] <= data_col54[32];
   data_col54[34] <= data_col54[33];
   data_col54[35] <= data_col54[34];
   data_col54[36] <= data_col54[35];
   data_col54[37] <= data_col54[36];
   data_col54[38] <= data_col54[37];
   data_col54[39] <= data_col54[38];
   data_col54[40] <= data_col54[39];
   data_col54[41] <= data_col54[40];
   data_col54[42] <= data_col54[41];
   data_col54[43] <= data_col54[42];
   data_col54[44] <= data_col54[43];
   data_col54[45] <= data_col54[44];
   data_col54[46] <= data_col54[45];
   data_col54[47] <= data_col54[46];
   data_col54[48] <= data_col54[47];
   data_col54[49] <= data_col54[48];
   data_col54[50] <= data_col54[49];
   data_col54[51] <= data_col54[50];
   data_col54[52] <= data_col54[51];
   data_col54[53] <= data_col54[52];
   data_col54[54] <= data_col54[53];

   data_col55[1] <= data[45];
   data_col55[2] <= data_col55[1];
   data_col55[3] <= data_col55[2];
   data_col55[4] <= data_col55[3];
   data_col55[5] <= data_col55[4];
   data_col55[6] <= data_col55[5];
   data_col55[7] <= data_col55[6];
   data_col55[8] <= data_col55[7];
   data_col55[9] <= data_col55[8];
   data_col55[10] <= data_col55[9];
   data_col55[11] <= data_col55[10];
   data_col55[12] <= data_col55[11];
   data_col55[13] <= data_col55[12];
   data_col55[14] <= data_col55[13];
   data_col55[15] <= data_col55[14];
   data_col55[16] <= data_col55[15];
   data_col55[17] <= data_col55[16];
   data_col55[18] <= data_col55[17];
   data_col55[19] <= data_col55[18];
   data_col55[20] <= data_col55[19];
   data_col55[21] <= data_col55[20];
   data_col55[22] <= data_col55[21];
   data_col55[23] <= data_col55[22];
   data_col55[24] <= data_col55[23];
   data_col55[25] <= data_col55[24];
   data_col55[26] <= data_col55[25];
   data_col55[27] <= data_col55[26];
   data_col55[28] <= data_col55[27];
   data_col55[29] <= data_col55[28];
   data_col55[30] <= data_col55[29];
   data_col55[31] <= data_col55[30];
   data_col55[32] <= data_col55[31];
   data_col55[33] <= data_col55[32];
   data_col55[34] <= data_col55[33];
   data_col55[35] <= data_col55[34];
   data_col55[36] <= data_col55[35];
   data_col55[37] <= data_col55[36];
   data_col55[38] <= data_col55[37];
   data_col55[39] <= data_col55[38];
   data_col55[40] <= data_col55[39];
   data_col55[41] <= data_col55[40];
   data_col55[42] <= data_col55[41];
   data_col55[43] <= data_col55[42];
   data_col55[44] <= data_col55[43];
   data_col55[45] <= data_col55[44];
   data_col55[46] <= data_col55[45];
   data_col55[47] <= data_col55[46];
   data_col55[48] <= data_col55[47];
   data_col55[49] <= data_col55[48];
   data_col55[50] <= data_col55[49];
   data_col55[51] <= data_col55[50];
   data_col55[52] <= data_col55[51];
   data_col55[53] <= data_col55[52];
   data_col55[54] <= data_col55[53];
   data_col55[55] <= data_col55[54];

   data_col56[1] <= data[44];
   data_col56[2] <= data_col56[1];
   data_col56[3] <= data_col56[2];
   data_col56[4] <= data_col56[3];
   data_col56[5] <= data_col56[4];
   data_col56[6] <= data_col56[5];
   data_col56[7] <= data_col56[6];
   data_col56[8] <= data_col56[7];
   data_col56[9] <= data_col56[8];
   data_col56[10] <= data_col56[9];
   data_col56[11] <= data_col56[10];
   data_col56[12] <= data_col56[11];
   data_col56[13] <= data_col56[12];
   data_col56[14] <= data_col56[13];
   data_col56[15] <= data_col56[14];
   data_col56[16] <= data_col56[15];
   data_col56[17] <= data_col56[16];
   data_col56[18] <= data_col56[17];
   data_col56[19] <= data_col56[18];
   data_col56[20] <= data_col56[19];
   data_col56[21] <= data_col56[20];
   data_col56[22] <= data_col56[21];
   data_col56[23] <= data_col56[22];
   data_col56[24] <= data_col56[23];
   data_col56[25] <= data_col56[24];
   data_col56[26] <= data_col56[25];
   data_col56[27] <= data_col56[26];
   data_col56[28] <= data_col56[27];
   data_col56[29] <= data_col56[28];
   data_col56[30] <= data_col56[29];
   data_col56[31] <= data_col56[30];
   data_col56[32] <= data_col56[31];
   data_col56[33] <= data_col56[32];
   data_col56[34] <= data_col56[33];
   data_col56[35] <= data_col56[34];
   data_col56[36] <= data_col56[35];
   data_col56[37] <= data_col56[36];
   data_col56[38] <= data_col56[37];
   data_col56[39] <= data_col56[38];
   data_col56[40] <= data_col56[39];
   data_col56[41] <= data_col56[40];
   data_col56[42] <= data_col56[41];
   data_col56[43] <= data_col56[42];
   data_col56[44] <= data_col56[43];
   data_col56[45] <= data_col56[44];
   data_col56[46] <= data_col56[45];
   data_col56[47] <= data_col56[46];
   data_col56[48] <= data_col56[47];
   data_col56[49] <= data_col56[48];
   data_col56[50] <= data_col56[49];
   data_col56[51] <= data_col56[50];
   data_col56[52] <= data_col56[51];
   data_col56[53] <= data_col56[52];
   data_col56[54] <= data_col56[53];
   data_col56[55] <= data_col56[54];
   data_col56[56] <= data_col56[55];

   data_col57[1] <= data[43];
   data_col57[2] <= data_col57[1];
   data_col57[3] <= data_col57[2];
   data_col57[4] <= data_col57[3];
   data_col57[5] <= data_col57[4];
   data_col57[6] <= data_col57[5];
   data_col57[7] <= data_col57[6];
   data_col57[8] <= data_col57[7];
   data_col57[9] <= data_col57[8];
   data_col57[10] <= data_col57[9];
   data_col57[11] <= data_col57[10];
   data_col57[12] <= data_col57[11];
   data_col57[13] <= data_col57[12];
   data_col57[14] <= data_col57[13];
   data_col57[15] <= data_col57[14];
   data_col57[16] <= data_col57[15];
   data_col57[17] <= data_col57[16];
   data_col57[18] <= data_col57[17];
   data_col57[19] <= data_col57[18];
   data_col57[20] <= data_col57[19];
   data_col57[21] <= data_col57[20];
   data_col57[22] <= data_col57[21];
   data_col57[23] <= data_col57[22];
   data_col57[24] <= data_col57[23];
   data_col57[25] <= data_col57[24];
   data_col57[26] <= data_col57[25];
   data_col57[27] <= data_col57[26];
   data_col57[28] <= data_col57[27];
   data_col57[29] <= data_col57[28];
   data_col57[30] <= data_col57[29];
   data_col57[31] <= data_col57[30];
   data_col57[32] <= data_col57[31];
   data_col57[33] <= data_col57[32];
   data_col57[34] <= data_col57[33];
   data_col57[35] <= data_col57[34];
   data_col57[36] <= data_col57[35];
   data_col57[37] <= data_col57[36];
   data_col57[38] <= data_col57[37];
   data_col57[39] <= data_col57[38];
   data_col57[40] <= data_col57[39];
   data_col57[41] <= data_col57[40];
   data_col57[42] <= data_col57[41];
   data_col57[43] <= data_col57[42];
   data_col57[44] <= data_col57[43];
   data_col57[45] <= data_col57[44];
   data_col57[46] <= data_col57[45];
   data_col57[47] <= data_col57[46];
   data_col57[48] <= data_col57[47];
   data_col57[49] <= data_col57[48];
   data_col57[50] <= data_col57[49];
   data_col57[51] <= data_col57[50];
   data_col57[52] <= data_col57[51];
   data_col57[53] <= data_col57[52];
   data_col57[54] <= data_col57[53];
   data_col57[55] <= data_col57[54];
   data_col57[56] <= data_col57[55];
   data_col57[57] <= data_col57[56];

   data_col58[1] <= data[42];
   data_col58[2] <= data_col58[1];
   data_col58[3] <= data_col58[2];
   data_col58[4] <= data_col58[3];
   data_col58[5] <= data_col58[4];
   data_col58[6] <= data_col58[5];
   data_col58[7] <= data_col58[6];
   data_col58[8] <= data_col58[7];
   data_col58[9] <= data_col58[8];
   data_col58[10] <= data_col58[9];
   data_col58[11] <= data_col58[10];
   data_col58[12] <= data_col58[11];
   data_col58[13] <= data_col58[12];
   data_col58[14] <= data_col58[13];
   data_col58[15] <= data_col58[14];
   data_col58[16] <= data_col58[15];
   data_col58[17] <= data_col58[16];
   data_col58[18] <= data_col58[17];
   data_col58[19] <= data_col58[18];
   data_col58[20] <= data_col58[19];
   data_col58[21] <= data_col58[20];
   data_col58[22] <= data_col58[21];
   data_col58[23] <= data_col58[22];
   data_col58[24] <= data_col58[23];
   data_col58[25] <= data_col58[24];
   data_col58[26] <= data_col58[25];
   data_col58[27] <= data_col58[26];
   data_col58[28] <= data_col58[27];
   data_col58[29] <= data_col58[28];
   data_col58[30] <= data_col58[29];
   data_col58[31] <= data_col58[30];
   data_col58[32] <= data_col58[31];
   data_col58[33] <= data_col58[32];
   data_col58[34] <= data_col58[33];
   data_col58[35] <= data_col58[34];
   data_col58[36] <= data_col58[35];
   data_col58[37] <= data_col58[36];
   data_col58[38] <= data_col58[37];
   data_col58[39] <= data_col58[38];
   data_col58[40] <= data_col58[39];
   data_col58[41] <= data_col58[40];
   data_col58[42] <= data_col58[41];
   data_col58[43] <= data_col58[42];
   data_col58[44] <= data_col58[43];
   data_col58[45] <= data_col58[44];
   data_col58[46] <= data_col58[45];
   data_col58[47] <= data_col58[46];
   data_col58[48] <= data_col58[47];
   data_col58[49] <= data_col58[48];
   data_col58[50] <= data_col58[49];
   data_col58[51] <= data_col58[50];
   data_col58[52] <= data_col58[51];
   data_col58[53] <= data_col58[52];
   data_col58[54] <= data_col58[53];
   data_col58[55] <= data_col58[54];
   data_col58[56] <= data_col58[55];
   data_col58[57] <= data_col58[56];
   data_col58[58] <= data_col58[57];

   data_col59[1] <= data[41];
   data_col59[2] <= data_col59[1];
   data_col59[3] <= data_col59[2];
   data_col59[4] <= data_col59[3];
   data_col59[5] <= data_col59[4];
   data_col59[6] <= data_col59[5];
   data_col59[7] <= data_col59[6];
   data_col59[8] <= data_col59[7];
   data_col59[9] <= data_col59[8];
   data_col59[10] <= data_col59[9];
   data_col59[11] <= data_col59[10];
   data_col59[12] <= data_col59[11];
   data_col59[13] <= data_col59[12];
   data_col59[14] <= data_col59[13];
   data_col59[15] <= data_col59[14];
   data_col59[16] <= data_col59[15];
   data_col59[17] <= data_col59[16];
   data_col59[18] <= data_col59[17];
   data_col59[19] <= data_col59[18];
   data_col59[20] <= data_col59[19];
   data_col59[21] <= data_col59[20];
   data_col59[22] <= data_col59[21];
   data_col59[23] <= data_col59[22];
   data_col59[24] <= data_col59[23];
   data_col59[25] <= data_col59[24];
   data_col59[26] <= data_col59[25];
   data_col59[27] <= data_col59[26];
   data_col59[28] <= data_col59[27];
   data_col59[29] <= data_col59[28];
   data_col59[30] <= data_col59[29];
   data_col59[31] <= data_col59[30];
   data_col59[32] <= data_col59[31];
   data_col59[33] <= data_col59[32];
   data_col59[34] <= data_col59[33];
   data_col59[35] <= data_col59[34];
   data_col59[36] <= data_col59[35];
   data_col59[37] <= data_col59[36];
   data_col59[38] <= data_col59[37];
   data_col59[39] <= data_col59[38];
   data_col59[40] <= data_col59[39];
   data_col59[41] <= data_col59[40];
   data_col59[42] <= data_col59[41];
   data_col59[43] <= data_col59[42];
   data_col59[44] <= data_col59[43];
   data_col59[45] <= data_col59[44];
   data_col59[46] <= data_col59[45];
   data_col59[47] <= data_col59[46];
   data_col59[48] <= data_col59[47];
   data_col59[49] <= data_col59[48];
   data_col59[50] <= data_col59[49];
   data_col59[51] <= data_col59[50];
   data_col59[52] <= data_col59[51];
   data_col59[53] <= data_col59[52];
   data_col59[54] <= data_col59[53];
   data_col59[55] <= data_col59[54];
   data_col59[56] <= data_col59[55];
   data_col59[57] <= data_col59[56];
   data_col59[58] <= data_col59[57];
   data_col59[59] <= data_col59[58];

   data_col60[1] <= data[40];
   data_col60[2] <= data_col60[1];
   data_col60[3] <= data_col60[2];
   data_col60[4] <= data_col60[3];
   data_col60[5] <= data_col60[4];
   data_col60[6] <= data_col60[5];
   data_col60[7] <= data_col60[6];
   data_col60[8] <= data_col60[7];
   data_col60[9] <= data_col60[8];
   data_col60[10] <= data_col60[9];
   data_col60[11] <= data_col60[10];
   data_col60[12] <= data_col60[11];
   data_col60[13] <= data_col60[12];
   data_col60[14] <= data_col60[13];
   data_col60[15] <= data_col60[14];
   data_col60[16] <= data_col60[15];
   data_col60[17] <= data_col60[16];
   data_col60[18] <= data_col60[17];
   data_col60[19] <= data_col60[18];
   data_col60[20] <= data_col60[19];
   data_col60[21] <= data_col60[20];
   data_col60[22] <= data_col60[21];
   data_col60[23] <= data_col60[22];
   data_col60[24] <= data_col60[23];
   data_col60[25] <= data_col60[24];
   data_col60[26] <= data_col60[25];
   data_col60[27] <= data_col60[26];
   data_col60[28] <= data_col60[27];
   data_col60[29] <= data_col60[28];
   data_col60[30] <= data_col60[29];
   data_col60[31] <= data_col60[30];
   data_col60[32] <= data_col60[31];
   data_col60[33] <= data_col60[32];
   data_col60[34] <= data_col60[33];
   data_col60[35] <= data_col60[34];
   data_col60[36] <= data_col60[35];
   data_col60[37] <= data_col60[36];
   data_col60[38] <= data_col60[37];
   data_col60[39] <= data_col60[38];
   data_col60[40] <= data_col60[39];
   data_col60[41] <= data_col60[40];
   data_col60[42] <= data_col60[41];
   data_col60[43] <= data_col60[42];
   data_col60[44] <= data_col60[43];
   data_col60[45] <= data_col60[44];
   data_col60[46] <= data_col60[45];
   data_col60[47] <= data_col60[46];
   data_col60[48] <= data_col60[47];
   data_col60[49] <= data_col60[48];
   data_col60[50] <= data_col60[49];
   data_col60[51] <= data_col60[50];
   data_col60[52] <= data_col60[51];
   data_col60[53] <= data_col60[52];
   data_col60[54] <= data_col60[53];
   data_col60[55] <= data_col60[54];
   data_col60[56] <= data_col60[55];
   data_col60[57] <= data_col60[56];
   data_col60[58] <= data_col60[57];
   data_col60[59] <= data_col60[58];
   data_col60[60] <= data_col60[59];

   data_col61[1] <= data[39];
   data_col61[2] <= data_col61[1];
   data_col61[3] <= data_col61[2];
   data_col61[4] <= data_col61[3];
   data_col61[5] <= data_col61[4];
   data_col61[6] <= data_col61[5];
   data_col61[7] <= data_col61[6];
   data_col61[8] <= data_col61[7];
   data_col61[9] <= data_col61[8];
   data_col61[10] <= data_col61[9];
   data_col61[11] <= data_col61[10];
   data_col61[12] <= data_col61[11];
   data_col61[13] <= data_col61[12];
   data_col61[14] <= data_col61[13];
   data_col61[15] <= data_col61[14];
   data_col61[16] <= data_col61[15];
   data_col61[17] <= data_col61[16];
   data_col61[18] <= data_col61[17];
   data_col61[19] <= data_col61[18];
   data_col61[20] <= data_col61[19];
   data_col61[21] <= data_col61[20];
   data_col61[22] <= data_col61[21];
   data_col61[23] <= data_col61[22];
   data_col61[24] <= data_col61[23];
   data_col61[25] <= data_col61[24];
   data_col61[26] <= data_col61[25];
   data_col61[27] <= data_col61[26];
   data_col61[28] <= data_col61[27];
   data_col61[29] <= data_col61[28];
   data_col61[30] <= data_col61[29];
   data_col61[31] <= data_col61[30];
   data_col61[32] <= data_col61[31];
   data_col61[33] <= data_col61[32];
   data_col61[34] <= data_col61[33];
   data_col61[35] <= data_col61[34];
   data_col61[36] <= data_col61[35];
   data_col61[37] <= data_col61[36];
   data_col61[38] <= data_col61[37];
   data_col61[39] <= data_col61[38];
   data_col61[40] <= data_col61[39];
   data_col61[41] <= data_col61[40];
   data_col61[42] <= data_col61[41];
   data_col61[43] <= data_col61[42];
   data_col61[44] <= data_col61[43];
   data_col61[45] <= data_col61[44];
   data_col61[46] <= data_col61[45];
   data_col61[47] <= data_col61[46];
   data_col61[48] <= data_col61[47];
   data_col61[49] <= data_col61[48];
   data_col61[50] <= data_col61[49];
   data_col61[51] <= data_col61[50];
   data_col61[52] <= data_col61[51];
   data_col61[53] <= data_col61[52];
   data_col61[54] <= data_col61[53];
   data_col61[55] <= data_col61[54];
   data_col61[56] <= data_col61[55];
   data_col61[57] <= data_col61[56];
   data_col61[58] <= data_col61[57];
   data_col61[59] <= data_col61[58];
   data_col61[60] <= data_col61[59];
   data_col61[61] <= data_col61[60];

   data_col62[1] <= data[38];
   data_col62[2] <= data_col62[1];
   data_col62[3] <= data_col62[2];
   data_col62[4] <= data_col62[3];
   data_col62[5] <= data_col62[4];
   data_col62[6] <= data_col62[5];
   data_col62[7] <= data_col62[6];
   data_col62[8] <= data_col62[7];
   data_col62[9] <= data_col62[8];
   data_col62[10] <= data_col62[9];
   data_col62[11] <= data_col62[10];
   data_col62[12] <= data_col62[11];
   data_col62[13] <= data_col62[12];
   data_col62[14] <= data_col62[13];
   data_col62[15] <= data_col62[14];
   data_col62[16] <= data_col62[15];
   data_col62[17] <= data_col62[16];
   data_col62[18] <= data_col62[17];
   data_col62[19] <= data_col62[18];
   data_col62[20] <= data_col62[19];
   data_col62[21] <= data_col62[20];
   data_col62[22] <= data_col62[21];
   data_col62[23] <= data_col62[22];
   data_col62[24] <= data_col62[23];
   data_col62[25] <= data_col62[24];
   data_col62[26] <= data_col62[25];
   data_col62[27] <= data_col62[26];
   data_col62[28] <= data_col62[27];
   data_col62[29] <= data_col62[28];
   data_col62[30] <= data_col62[29];
   data_col62[31] <= data_col62[30];
   data_col62[32] <= data_col62[31];
   data_col62[33] <= data_col62[32];
   data_col62[34] <= data_col62[33];
   data_col62[35] <= data_col62[34];
   data_col62[36] <= data_col62[35];
   data_col62[37] <= data_col62[36];
   data_col62[38] <= data_col62[37];
   data_col62[39] <= data_col62[38];
   data_col62[40] <= data_col62[39];
   data_col62[41] <= data_col62[40];
   data_col62[42] <= data_col62[41];
   data_col62[43] <= data_col62[42];
   data_col62[44] <= data_col62[43];
   data_col62[45] <= data_col62[44];
   data_col62[46] <= data_col62[45];
   data_col62[47] <= data_col62[46];
   data_col62[48] <= data_col62[47];
   data_col62[49] <= data_col62[48];
   data_col62[50] <= data_col62[49];
   data_col62[51] <= data_col62[50];
   data_col62[52] <= data_col62[51];
   data_col62[53] <= data_col62[52];
   data_col62[54] <= data_col62[53];
   data_col62[55] <= data_col62[54];
   data_col62[56] <= data_col62[55];
   data_col62[57] <= data_col62[56];
   data_col62[58] <= data_col62[57];
   data_col62[59] <= data_col62[58];
   data_col62[60] <= data_col62[59];
   data_col62[61] <= data_col62[60];
   data_col62[62] <= data_col62[61];

   data_col63[1] <= data[37];
   data_col63[2] <= data_col63[1];
   data_col63[3] <= data_col63[2];
   data_col63[4] <= data_col63[3];
   data_col63[5] <= data_col63[4];
   data_col63[6] <= data_col63[5];
   data_col63[7] <= data_col63[6];
   data_col63[8] <= data_col63[7];
   data_col63[9] <= data_col63[8];
   data_col63[10] <= data_col63[9];
   data_col63[11] <= data_col63[10];
   data_col63[12] <= data_col63[11];
   data_col63[13] <= data_col63[12];
   data_col63[14] <= data_col63[13];
   data_col63[15] <= data_col63[14];
   data_col63[16] <= data_col63[15];
   data_col63[17] <= data_col63[16];
   data_col63[18] <= data_col63[17];
   data_col63[19] <= data_col63[18];
   data_col63[20] <= data_col63[19];
   data_col63[21] <= data_col63[20];
   data_col63[22] <= data_col63[21];
   data_col63[23] <= data_col63[22];
   data_col63[24] <= data_col63[23];
   data_col63[25] <= data_col63[24];
   data_col63[26] <= data_col63[25];
   data_col63[27] <= data_col63[26];
   data_col63[28] <= data_col63[27];
   data_col63[29] <= data_col63[28];
   data_col63[30] <= data_col63[29];
   data_col63[31] <= data_col63[30];
   data_col63[32] <= data_col63[31];
   data_col63[33] <= data_col63[32];
   data_col63[34] <= data_col63[33];
   data_col63[35] <= data_col63[34];
   data_col63[36] <= data_col63[35];
   data_col63[37] <= data_col63[36];
   data_col63[38] <= data_col63[37];
   data_col63[39] <= data_col63[38];
   data_col63[40] <= data_col63[39];
   data_col63[41] <= data_col63[40];
   data_col63[42] <= data_col63[41];
   data_col63[43] <= data_col63[42];
   data_col63[44] <= data_col63[43];
   data_col63[45] <= data_col63[44];
   data_col63[46] <= data_col63[45];
   data_col63[47] <= data_col63[46];
   data_col63[48] <= data_col63[47];
   data_col63[49] <= data_col63[48];
   data_col63[50] <= data_col63[49];
   data_col63[51] <= data_col63[50];
   data_col63[52] <= data_col63[51];
   data_col63[53] <= data_col63[52];
   data_col63[54] <= data_col63[53];
   data_col63[55] <= data_col63[54];
   data_col63[56] <= data_col63[55];
   data_col63[57] <= data_col63[56];
   data_col63[58] <= data_col63[57];
   data_col63[59] <= data_col63[58];
   data_col63[60] <= data_col63[59];
   data_col63[61] <= data_col63[60];
   data_col63[62] <= data_col63[61];
   data_col63[63] <= data_col63[62];

   data_col64[1] <= data[36];
   data_col64[2] <= data_col64[1];
   data_col64[3] <= data_col64[2];
   data_col64[4] <= data_col64[3];
   data_col64[5] <= data_col64[4];
   data_col64[6] <= data_col64[5];
   data_col64[7] <= data_col64[6];
   data_col64[8] <= data_col64[7];
   data_col64[9] <= data_col64[8];
   data_col64[10] <= data_col64[9];
   data_col64[11] <= data_col64[10];
   data_col64[12] <= data_col64[11];
   data_col64[13] <= data_col64[12];
   data_col64[14] <= data_col64[13];
   data_col64[15] <= data_col64[14];
   data_col64[16] <= data_col64[15];
   data_col64[17] <= data_col64[16];
   data_col64[18] <= data_col64[17];
   data_col64[19] <= data_col64[18];
   data_col64[20] <= data_col64[19];
   data_col64[21] <= data_col64[20];
   data_col64[22] <= data_col64[21];
   data_col64[23] <= data_col64[22];
   data_col64[24] <= data_col64[23];
   data_col64[25] <= data_col64[24];
   data_col64[26] <= data_col64[25];
   data_col64[27] <= data_col64[26];
   data_col64[28] <= data_col64[27];
   data_col64[29] <= data_col64[28];
   data_col64[30] <= data_col64[29];
   data_col64[31] <= data_col64[30];
   data_col64[32] <= data_col64[31];
   data_col64[33] <= data_col64[32];
   data_col64[34] <= data_col64[33];
   data_col64[35] <= data_col64[34];
   data_col64[36] <= data_col64[35];
   data_col64[37] <= data_col64[36];
   data_col64[38] <= data_col64[37];
   data_col64[39] <= data_col64[38];
   data_col64[40] <= data_col64[39];
   data_col64[41] <= data_col64[40];
   data_col64[42] <= data_col64[41];
   data_col64[43] <= data_col64[42];
   data_col64[44] <= data_col64[43];
   data_col64[45] <= data_col64[44];
   data_col64[46] <= data_col64[45];
   data_col64[47] <= data_col64[46];
   data_col64[48] <= data_col64[47];
   data_col64[49] <= data_col64[48];
   data_col64[50] <= data_col64[49];
   data_col64[51] <= data_col64[50];
   data_col64[52] <= data_col64[51];
   data_col64[53] <= data_col64[52];
   data_col64[54] <= data_col64[53];
   data_col64[55] <= data_col64[54];
   data_col64[56] <= data_col64[55];
   data_col64[57] <= data_col64[56];
   data_col64[58] <= data_col64[57];
   data_col64[59] <= data_col64[58];
   data_col64[60] <= data_col64[59];
   data_col64[61] <= data_col64[60];
   data_col64[62] <= data_col64[61];
   data_col64[63] <= data_col64[62];
   data_col64[64] <= data_col64[63];

   data_col65[1] <= data[35];
   data_col65[2] <= data_col65[1];
   data_col65[3] <= data_col65[2];
   data_col65[4] <= data_col65[3];
   data_col65[5] <= data_col65[4];
   data_col65[6] <= data_col65[5];
   data_col65[7] <= data_col65[6];
   data_col65[8] <= data_col65[7];
   data_col65[9] <= data_col65[8];
   data_col65[10] <= data_col65[9];
   data_col65[11] <= data_col65[10];
   data_col65[12] <= data_col65[11];
   data_col65[13] <= data_col65[12];
   data_col65[14] <= data_col65[13];
   data_col65[15] <= data_col65[14];
   data_col65[16] <= data_col65[15];
   data_col65[17] <= data_col65[16];
   data_col65[18] <= data_col65[17];
   data_col65[19] <= data_col65[18];
   data_col65[20] <= data_col65[19];
   data_col65[21] <= data_col65[20];
   data_col65[22] <= data_col65[21];
   data_col65[23] <= data_col65[22];
   data_col65[24] <= data_col65[23];
   data_col65[25] <= data_col65[24];
   data_col65[26] <= data_col65[25];
   data_col65[27] <= data_col65[26];
   data_col65[28] <= data_col65[27];
   data_col65[29] <= data_col65[28];
   data_col65[30] <= data_col65[29];
   data_col65[31] <= data_col65[30];
   data_col65[32] <= data_col65[31];
   data_col65[33] <= data_col65[32];
   data_col65[34] <= data_col65[33];
   data_col65[35] <= data_col65[34];
   data_col65[36] <= data_col65[35];
   data_col65[37] <= data_col65[36];
   data_col65[38] <= data_col65[37];
   data_col65[39] <= data_col65[38];
   data_col65[40] <= data_col65[39];
   data_col65[41] <= data_col65[40];
   data_col65[42] <= data_col65[41];
   data_col65[43] <= data_col65[42];
   data_col65[44] <= data_col65[43];
   data_col65[45] <= data_col65[44];
   data_col65[46] <= data_col65[45];
   data_col65[47] <= data_col65[46];
   data_col65[48] <= data_col65[47];
   data_col65[49] <= data_col65[48];
   data_col65[50] <= data_col65[49];
   data_col65[51] <= data_col65[50];
   data_col65[52] <= data_col65[51];
   data_col65[53] <= data_col65[52];
   data_col65[54] <= data_col65[53];
   data_col65[55] <= data_col65[54];
   data_col65[56] <= data_col65[55];
   data_col65[57] <= data_col65[56];
   data_col65[58] <= data_col65[57];
   data_col65[59] <= data_col65[58];
   data_col65[60] <= data_col65[59];
   data_col65[61] <= data_col65[60];
   data_col65[62] <= data_col65[61];
   data_col65[63] <= data_col65[62];
   data_col65[64] <= data_col65[63];
   data_col65[65] <= data_col65[64];

   data_col66[1] <= data[34];
   data_col66[2] <= data_col66[1];
   data_col66[3] <= data_col66[2];
   data_col66[4] <= data_col66[3];
   data_col66[5] <= data_col66[4];
   data_col66[6] <= data_col66[5];
   data_col66[7] <= data_col66[6];
   data_col66[8] <= data_col66[7];
   data_col66[9] <= data_col66[8];
   data_col66[10] <= data_col66[9];
   data_col66[11] <= data_col66[10];
   data_col66[12] <= data_col66[11];
   data_col66[13] <= data_col66[12];
   data_col66[14] <= data_col66[13];
   data_col66[15] <= data_col66[14];
   data_col66[16] <= data_col66[15];
   data_col66[17] <= data_col66[16];
   data_col66[18] <= data_col66[17];
   data_col66[19] <= data_col66[18];
   data_col66[20] <= data_col66[19];
   data_col66[21] <= data_col66[20];
   data_col66[22] <= data_col66[21];
   data_col66[23] <= data_col66[22];
   data_col66[24] <= data_col66[23];
   data_col66[25] <= data_col66[24];
   data_col66[26] <= data_col66[25];
   data_col66[27] <= data_col66[26];
   data_col66[28] <= data_col66[27];
   data_col66[29] <= data_col66[28];
   data_col66[30] <= data_col66[29];
   data_col66[31] <= data_col66[30];
   data_col66[32] <= data_col66[31];
   data_col66[33] <= data_col66[32];
   data_col66[34] <= data_col66[33];
   data_col66[35] <= data_col66[34];
   data_col66[36] <= data_col66[35];
   data_col66[37] <= data_col66[36];
   data_col66[38] <= data_col66[37];
   data_col66[39] <= data_col66[38];
   data_col66[40] <= data_col66[39];
   data_col66[41] <= data_col66[40];
   data_col66[42] <= data_col66[41];
   data_col66[43] <= data_col66[42];
   data_col66[44] <= data_col66[43];
   data_col66[45] <= data_col66[44];
   data_col66[46] <= data_col66[45];
   data_col66[47] <= data_col66[46];
   data_col66[48] <= data_col66[47];
   data_col66[49] <= data_col66[48];
   data_col66[50] <= data_col66[49];
   data_col66[51] <= data_col66[50];
   data_col66[52] <= data_col66[51];
   data_col66[53] <= data_col66[52];
   data_col66[54] <= data_col66[53];
   data_col66[55] <= data_col66[54];
   data_col66[56] <= data_col66[55];
   data_col66[57] <= data_col66[56];
   data_col66[58] <= data_col66[57];
   data_col66[59] <= data_col66[58];
   data_col66[60] <= data_col66[59];
   data_col66[61] <= data_col66[60];
   data_col66[62] <= data_col66[61];
   data_col66[63] <= data_col66[62];
   data_col66[64] <= data_col66[63];
   data_col66[65] <= data_col66[64];
   data_col66[66] <= data_col66[65];

   data_col67[1] <= data[33];
   data_col67[2] <= data_col67[1];
   data_col67[3] <= data_col67[2];
   data_col67[4] <= data_col67[3];
   data_col67[5] <= data_col67[4];
   data_col67[6] <= data_col67[5];
   data_col67[7] <= data_col67[6];
   data_col67[8] <= data_col67[7];
   data_col67[9] <= data_col67[8];
   data_col67[10] <= data_col67[9];
   data_col67[11] <= data_col67[10];
   data_col67[12] <= data_col67[11];
   data_col67[13] <= data_col67[12];
   data_col67[14] <= data_col67[13];
   data_col67[15] <= data_col67[14];
   data_col67[16] <= data_col67[15];
   data_col67[17] <= data_col67[16];
   data_col67[18] <= data_col67[17];
   data_col67[19] <= data_col67[18];
   data_col67[20] <= data_col67[19];
   data_col67[21] <= data_col67[20];
   data_col67[22] <= data_col67[21];
   data_col67[23] <= data_col67[22];
   data_col67[24] <= data_col67[23];
   data_col67[25] <= data_col67[24];
   data_col67[26] <= data_col67[25];
   data_col67[27] <= data_col67[26];
   data_col67[28] <= data_col67[27];
   data_col67[29] <= data_col67[28];
   data_col67[30] <= data_col67[29];
   data_col67[31] <= data_col67[30];
   data_col67[32] <= data_col67[31];
   data_col67[33] <= data_col67[32];
   data_col67[34] <= data_col67[33];
   data_col67[35] <= data_col67[34];
   data_col67[36] <= data_col67[35];
   data_col67[37] <= data_col67[36];
   data_col67[38] <= data_col67[37];
   data_col67[39] <= data_col67[38];
   data_col67[40] <= data_col67[39];
   data_col67[41] <= data_col67[40];
   data_col67[42] <= data_col67[41];
   data_col67[43] <= data_col67[42];
   data_col67[44] <= data_col67[43];
   data_col67[45] <= data_col67[44];
   data_col67[46] <= data_col67[45];
   data_col67[47] <= data_col67[46];
   data_col67[48] <= data_col67[47];
   data_col67[49] <= data_col67[48];
   data_col67[50] <= data_col67[49];
   data_col67[51] <= data_col67[50];
   data_col67[52] <= data_col67[51];
   data_col67[53] <= data_col67[52];
   data_col67[54] <= data_col67[53];
   data_col67[55] <= data_col67[54];
   data_col67[56] <= data_col67[55];
   data_col67[57] <= data_col67[56];
   data_col67[58] <= data_col67[57];
   data_col67[59] <= data_col67[58];
   data_col67[60] <= data_col67[59];
   data_col67[61] <= data_col67[60];
   data_col67[62] <= data_col67[61];
   data_col67[63] <= data_col67[62];
   data_col67[64] <= data_col67[63];
   data_col67[65] <= data_col67[64];
   data_col67[66] <= data_col67[65];
   data_col67[67] <= data_col67[66];

   data_col68[1] <= data[32];
   data_col68[2] <= data_col68[1];
   data_col68[3] <= data_col68[2];
   data_col68[4] <= data_col68[3];
   data_col68[5] <= data_col68[4];
   data_col68[6] <= data_col68[5];
   data_col68[7] <= data_col68[6];
   data_col68[8] <= data_col68[7];
   data_col68[9] <= data_col68[8];
   data_col68[10] <= data_col68[9];
   data_col68[11] <= data_col68[10];
   data_col68[12] <= data_col68[11];
   data_col68[13] <= data_col68[12];
   data_col68[14] <= data_col68[13];
   data_col68[15] <= data_col68[14];
   data_col68[16] <= data_col68[15];
   data_col68[17] <= data_col68[16];
   data_col68[18] <= data_col68[17];
   data_col68[19] <= data_col68[18];
   data_col68[20] <= data_col68[19];
   data_col68[21] <= data_col68[20];
   data_col68[22] <= data_col68[21];
   data_col68[23] <= data_col68[22];
   data_col68[24] <= data_col68[23];
   data_col68[25] <= data_col68[24];
   data_col68[26] <= data_col68[25];
   data_col68[27] <= data_col68[26];
   data_col68[28] <= data_col68[27];
   data_col68[29] <= data_col68[28];
   data_col68[30] <= data_col68[29];
   data_col68[31] <= data_col68[30];
   data_col68[32] <= data_col68[31];
   data_col68[33] <= data_col68[32];
   data_col68[34] <= data_col68[33];
   data_col68[35] <= data_col68[34];
   data_col68[36] <= data_col68[35];
   data_col68[37] <= data_col68[36];
   data_col68[38] <= data_col68[37];
   data_col68[39] <= data_col68[38];
   data_col68[40] <= data_col68[39];
   data_col68[41] <= data_col68[40];
   data_col68[42] <= data_col68[41];
   data_col68[43] <= data_col68[42];
   data_col68[44] <= data_col68[43];
   data_col68[45] <= data_col68[44];
   data_col68[46] <= data_col68[45];
   data_col68[47] <= data_col68[46];
   data_col68[48] <= data_col68[47];
   data_col68[49] <= data_col68[48];
   data_col68[50] <= data_col68[49];
   data_col68[51] <= data_col68[50];
   data_col68[52] <= data_col68[51];
   data_col68[53] <= data_col68[52];
   data_col68[54] <= data_col68[53];
   data_col68[55] <= data_col68[54];
   data_col68[56] <= data_col68[55];
   data_col68[57] <= data_col68[56];
   data_col68[58] <= data_col68[57];
   data_col68[59] <= data_col68[58];
   data_col68[60] <= data_col68[59];
   data_col68[61] <= data_col68[60];
   data_col68[62] <= data_col68[61];
   data_col68[63] <= data_col68[62];
   data_col68[64] <= data_col68[63];
   data_col68[65] <= data_col68[64];
   data_col68[66] <= data_col68[65];
   data_col68[67] <= data_col68[66];
   data_col68[68] <= data_col68[67];

   data_col69[1] <= data[31];
   data_col69[2] <= data_col69[1];
   data_col69[3] <= data_col69[2];
   data_col69[4] <= data_col69[3];
   data_col69[5] <= data_col69[4];
   data_col69[6] <= data_col69[5];
   data_col69[7] <= data_col69[6];
   data_col69[8] <= data_col69[7];
   data_col69[9] <= data_col69[8];
   data_col69[10] <= data_col69[9];
   data_col69[11] <= data_col69[10];
   data_col69[12] <= data_col69[11];
   data_col69[13] <= data_col69[12];
   data_col69[14] <= data_col69[13];
   data_col69[15] <= data_col69[14];
   data_col69[16] <= data_col69[15];
   data_col69[17] <= data_col69[16];
   data_col69[18] <= data_col69[17];
   data_col69[19] <= data_col69[18];
   data_col69[20] <= data_col69[19];
   data_col69[21] <= data_col69[20];
   data_col69[22] <= data_col69[21];
   data_col69[23] <= data_col69[22];
   data_col69[24] <= data_col69[23];
   data_col69[25] <= data_col69[24];
   data_col69[26] <= data_col69[25];
   data_col69[27] <= data_col69[26];
   data_col69[28] <= data_col69[27];
   data_col69[29] <= data_col69[28];
   data_col69[30] <= data_col69[29];
   data_col69[31] <= data_col69[30];
   data_col69[32] <= data_col69[31];
   data_col69[33] <= data_col69[32];
   data_col69[34] <= data_col69[33];
   data_col69[35] <= data_col69[34];
   data_col69[36] <= data_col69[35];
   data_col69[37] <= data_col69[36];
   data_col69[38] <= data_col69[37];
   data_col69[39] <= data_col69[38];
   data_col69[40] <= data_col69[39];
   data_col69[41] <= data_col69[40];
   data_col69[42] <= data_col69[41];
   data_col69[43] <= data_col69[42];
   data_col69[44] <= data_col69[43];
   data_col69[45] <= data_col69[44];
   data_col69[46] <= data_col69[45];
   data_col69[47] <= data_col69[46];
   data_col69[48] <= data_col69[47];
   data_col69[49] <= data_col69[48];
   data_col69[50] <= data_col69[49];
   data_col69[51] <= data_col69[50];
   data_col69[52] <= data_col69[51];
   data_col69[53] <= data_col69[52];
   data_col69[54] <= data_col69[53];
   data_col69[55] <= data_col69[54];
   data_col69[56] <= data_col69[55];
   data_col69[57] <= data_col69[56];
   data_col69[58] <= data_col69[57];
   data_col69[59] <= data_col69[58];
   data_col69[60] <= data_col69[59];
   data_col69[61] <= data_col69[60];
   data_col69[62] <= data_col69[61];
   data_col69[63] <= data_col69[62];
   data_col69[64] <= data_col69[63];
   data_col69[65] <= data_col69[64];
   data_col69[66] <= data_col69[65];
   data_col69[67] <= data_col69[66];
   data_col69[68] <= data_col69[67];
   data_col69[69] <= data_col69[68];

   data_col70[1] <= data[30];
   data_col70[2] <= data_col70[1];
   data_col70[3] <= data_col70[2];
   data_col70[4] <= data_col70[3];
   data_col70[5] <= data_col70[4];
   data_col70[6] <= data_col70[5];
   data_col70[7] <= data_col70[6];
   data_col70[8] <= data_col70[7];
   data_col70[9] <= data_col70[8];
   data_col70[10] <= data_col70[9];
   data_col70[11] <= data_col70[10];
   data_col70[12] <= data_col70[11];
   data_col70[13] <= data_col70[12];
   data_col70[14] <= data_col70[13];
   data_col70[15] <= data_col70[14];
   data_col70[16] <= data_col70[15];
   data_col70[17] <= data_col70[16];
   data_col70[18] <= data_col70[17];
   data_col70[19] <= data_col70[18];
   data_col70[20] <= data_col70[19];
   data_col70[21] <= data_col70[20];
   data_col70[22] <= data_col70[21];
   data_col70[23] <= data_col70[22];
   data_col70[24] <= data_col70[23];
   data_col70[25] <= data_col70[24];
   data_col70[26] <= data_col70[25];
   data_col70[27] <= data_col70[26];
   data_col70[28] <= data_col70[27];
   data_col70[29] <= data_col70[28];
   data_col70[30] <= data_col70[29];
   data_col70[31] <= data_col70[30];
   data_col70[32] <= data_col70[31];
   data_col70[33] <= data_col70[32];
   data_col70[34] <= data_col70[33];
   data_col70[35] <= data_col70[34];
   data_col70[36] <= data_col70[35];
   data_col70[37] <= data_col70[36];
   data_col70[38] <= data_col70[37];
   data_col70[39] <= data_col70[38];
   data_col70[40] <= data_col70[39];
   data_col70[41] <= data_col70[40];
   data_col70[42] <= data_col70[41];
   data_col70[43] <= data_col70[42];
   data_col70[44] <= data_col70[43];
   data_col70[45] <= data_col70[44];
   data_col70[46] <= data_col70[45];
   data_col70[47] <= data_col70[46];
   data_col70[48] <= data_col70[47];
   data_col70[49] <= data_col70[48];
   data_col70[50] <= data_col70[49];
   data_col70[51] <= data_col70[50];
   data_col70[52] <= data_col70[51];
   data_col70[53] <= data_col70[52];
   data_col70[54] <= data_col70[53];
   data_col70[55] <= data_col70[54];
   data_col70[56] <= data_col70[55];
   data_col70[57] <= data_col70[56];
   data_col70[58] <= data_col70[57];
   data_col70[59] <= data_col70[58];
   data_col70[60] <= data_col70[59];
   data_col70[61] <= data_col70[60];
   data_col70[62] <= data_col70[61];
   data_col70[63] <= data_col70[62];
   data_col70[64] <= data_col70[63];
   data_col70[65] <= data_col70[64];
   data_col70[66] <= data_col70[65];
   data_col70[67] <= data_col70[66];
   data_col70[68] <= data_col70[67];
   data_col70[69] <= data_col70[68];
   data_col70[70] <= data_col70[69];

   data_col71[1] <= data[29];
   data_col71[2] <= data_col71[1];
   data_col71[3] <= data_col71[2];
   data_col71[4] <= data_col71[3];
   data_col71[5] <= data_col71[4];
   data_col71[6] <= data_col71[5];
   data_col71[7] <= data_col71[6];
   data_col71[8] <= data_col71[7];
   data_col71[9] <= data_col71[8];
   data_col71[10] <= data_col71[9];
   data_col71[11] <= data_col71[10];
   data_col71[12] <= data_col71[11];
   data_col71[13] <= data_col71[12];
   data_col71[14] <= data_col71[13];
   data_col71[15] <= data_col71[14];
   data_col71[16] <= data_col71[15];
   data_col71[17] <= data_col71[16];
   data_col71[18] <= data_col71[17];
   data_col71[19] <= data_col71[18];
   data_col71[20] <= data_col71[19];
   data_col71[21] <= data_col71[20];
   data_col71[22] <= data_col71[21];
   data_col71[23] <= data_col71[22];
   data_col71[24] <= data_col71[23];
   data_col71[25] <= data_col71[24];
   data_col71[26] <= data_col71[25];
   data_col71[27] <= data_col71[26];
   data_col71[28] <= data_col71[27];
   data_col71[29] <= data_col71[28];
   data_col71[30] <= data_col71[29];
   data_col71[31] <= data_col71[30];
   data_col71[32] <= data_col71[31];
   data_col71[33] <= data_col71[32];
   data_col71[34] <= data_col71[33];
   data_col71[35] <= data_col71[34];
   data_col71[36] <= data_col71[35];
   data_col71[37] <= data_col71[36];
   data_col71[38] <= data_col71[37];
   data_col71[39] <= data_col71[38];
   data_col71[40] <= data_col71[39];
   data_col71[41] <= data_col71[40];
   data_col71[42] <= data_col71[41];
   data_col71[43] <= data_col71[42];
   data_col71[44] <= data_col71[43];
   data_col71[45] <= data_col71[44];
   data_col71[46] <= data_col71[45];
   data_col71[47] <= data_col71[46];
   data_col71[48] <= data_col71[47];
   data_col71[49] <= data_col71[48];
   data_col71[50] <= data_col71[49];
   data_col71[51] <= data_col71[50];
   data_col71[52] <= data_col71[51];
   data_col71[53] <= data_col71[52];
   data_col71[54] <= data_col71[53];
   data_col71[55] <= data_col71[54];
   data_col71[56] <= data_col71[55];
   data_col71[57] <= data_col71[56];
   data_col71[58] <= data_col71[57];
   data_col71[59] <= data_col71[58];
   data_col71[60] <= data_col71[59];
   data_col71[61] <= data_col71[60];
   data_col71[62] <= data_col71[61];
   data_col71[63] <= data_col71[62];
   data_col71[64] <= data_col71[63];
   data_col71[65] <= data_col71[64];
   data_col71[66] <= data_col71[65];
   data_col71[67] <= data_col71[66];
   data_col71[68] <= data_col71[67];
   data_col71[69] <= data_col71[68];
   data_col71[70] <= data_col71[69];
   data_col71[71] <= data_col71[70];

   data_col72[1] <= data[28];
   data_col72[2] <= data_col72[1];
   data_col72[3] <= data_col72[2];
   data_col72[4] <= data_col72[3];
   data_col72[5] <= data_col72[4];
   data_col72[6] <= data_col72[5];
   data_col72[7] <= data_col72[6];
   data_col72[8] <= data_col72[7];
   data_col72[9] <= data_col72[8];
   data_col72[10] <= data_col72[9];
   data_col72[11] <= data_col72[10];
   data_col72[12] <= data_col72[11];
   data_col72[13] <= data_col72[12];
   data_col72[14] <= data_col72[13];
   data_col72[15] <= data_col72[14];
   data_col72[16] <= data_col72[15];
   data_col72[17] <= data_col72[16];
   data_col72[18] <= data_col72[17];
   data_col72[19] <= data_col72[18];
   data_col72[20] <= data_col72[19];
   data_col72[21] <= data_col72[20];
   data_col72[22] <= data_col72[21];
   data_col72[23] <= data_col72[22];
   data_col72[24] <= data_col72[23];
   data_col72[25] <= data_col72[24];
   data_col72[26] <= data_col72[25];
   data_col72[27] <= data_col72[26];
   data_col72[28] <= data_col72[27];
   data_col72[29] <= data_col72[28];
   data_col72[30] <= data_col72[29];
   data_col72[31] <= data_col72[30];
   data_col72[32] <= data_col72[31];
   data_col72[33] <= data_col72[32];
   data_col72[34] <= data_col72[33];
   data_col72[35] <= data_col72[34];
   data_col72[36] <= data_col72[35];
   data_col72[37] <= data_col72[36];
   data_col72[38] <= data_col72[37];
   data_col72[39] <= data_col72[38];
   data_col72[40] <= data_col72[39];
   data_col72[41] <= data_col72[40];
   data_col72[42] <= data_col72[41];
   data_col72[43] <= data_col72[42];
   data_col72[44] <= data_col72[43];
   data_col72[45] <= data_col72[44];
   data_col72[46] <= data_col72[45];
   data_col72[47] <= data_col72[46];
   data_col72[48] <= data_col72[47];
   data_col72[49] <= data_col72[48];
   data_col72[50] <= data_col72[49];
   data_col72[51] <= data_col72[50];
   data_col72[52] <= data_col72[51];
   data_col72[53] <= data_col72[52];
   data_col72[54] <= data_col72[53];
   data_col72[55] <= data_col72[54];
   data_col72[56] <= data_col72[55];
   data_col72[57] <= data_col72[56];
   data_col72[58] <= data_col72[57];
   data_col72[59] <= data_col72[58];
   data_col72[60] <= data_col72[59];
   data_col72[61] <= data_col72[60];
   data_col72[62] <= data_col72[61];
   data_col72[63] <= data_col72[62];
   data_col72[64] <= data_col72[63];
   data_col72[65] <= data_col72[64];
   data_col72[66] <= data_col72[65];
   data_col72[67] <= data_col72[66];
   data_col72[68] <= data_col72[67];
   data_col72[69] <= data_col72[68];
   data_col72[70] <= data_col72[69];
   data_col72[71] <= data_col72[70];
   data_col72[72] <= data_col72[71];

   data_col73[1] <= data[27];
   data_col73[2] <= data_col73[1];
   data_col73[3] <= data_col73[2];
   data_col73[4] <= data_col73[3];
   data_col73[5] <= data_col73[4];
   data_col73[6] <= data_col73[5];
   data_col73[7] <= data_col73[6];
   data_col73[8] <= data_col73[7];
   data_col73[9] <= data_col73[8];
   data_col73[10] <= data_col73[9];
   data_col73[11] <= data_col73[10];
   data_col73[12] <= data_col73[11];
   data_col73[13] <= data_col73[12];
   data_col73[14] <= data_col73[13];
   data_col73[15] <= data_col73[14];
   data_col73[16] <= data_col73[15];
   data_col73[17] <= data_col73[16];
   data_col73[18] <= data_col73[17];
   data_col73[19] <= data_col73[18];
   data_col73[20] <= data_col73[19];
   data_col73[21] <= data_col73[20];
   data_col73[22] <= data_col73[21];
   data_col73[23] <= data_col73[22];
   data_col73[24] <= data_col73[23];
   data_col73[25] <= data_col73[24];
   data_col73[26] <= data_col73[25];
   data_col73[27] <= data_col73[26];
   data_col73[28] <= data_col73[27];
   data_col73[29] <= data_col73[28];
   data_col73[30] <= data_col73[29];
   data_col73[31] <= data_col73[30];
   data_col73[32] <= data_col73[31];
   data_col73[33] <= data_col73[32];
   data_col73[34] <= data_col73[33];
   data_col73[35] <= data_col73[34];
   data_col73[36] <= data_col73[35];
   data_col73[37] <= data_col73[36];
   data_col73[38] <= data_col73[37];
   data_col73[39] <= data_col73[38];
   data_col73[40] <= data_col73[39];
   data_col73[41] <= data_col73[40];
   data_col73[42] <= data_col73[41];
   data_col73[43] <= data_col73[42];
   data_col73[44] <= data_col73[43];
   data_col73[45] <= data_col73[44];
   data_col73[46] <= data_col73[45];
   data_col73[47] <= data_col73[46];
   data_col73[48] <= data_col73[47];
   data_col73[49] <= data_col73[48];
   data_col73[50] <= data_col73[49];
   data_col73[51] <= data_col73[50];
   data_col73[52] <= data_col73[51];
   data_col73[53] <= data_col73[52];
   data_col73[54] <= data_col73[53];
   data_col73[55] <= data_col73[54];
   data_col73[56] <= data_col73[55];
   data_col73[57] <= data_col73[56];
   data_col73[58] <= data_col73[57];
   data_col73[59] <= data_col73[58];
   data_col73[60] <= data_col73[59];
   data_col73[61] <= data_col73[60];
   data_col73[62] <= data_col73[61];
   data_col73[63] <= data_col73[62];
   data_col73[64] <= data_col73[63];
   data_col73[65] <= data_col73[64];
   data_col73[66] <= data_col73[65];
   data_col73[67] <= data_col73[66];
   data_col73[68] <= data_col73[67];
   data_col73[69] <= data_col73[68];
   data_col73[70] <= data_col73[69];
   data_col73[71] <= data_col73[70];
   data_col73[72] <= data_col73[71];
   data_col73[73] <= data_col73[72];

   data_col74[1] <= data[26];
   data_col74[2] <= data_col74[1];
   data_col74[3] <= data_col74[2];
   data_col74[4] <= data_col74[3];
   data_col74[5] <= data_col74[4];
   data_col74[6] <= data_col74[5];
   data_col74[7] <= data_col74[6];
   data_col74[8] <= data_col74[7];
   data_col74[9] <= data_col74[8];
   data_col74[10] <= data_col74[9];
   data_col74[11] <= data_col74[10];
   data_col74[12] <= data_col74[11];
   data_col74[13] <= data_col74[12];
   data_col74[14] <= data_col74[13];
   data_col74[15] <= data_col74[14];
   data_col74[16] <= data_col74[15];
   data_col74[17] <= data_col74[16];
   data_col74[18] <= data_col74[17];
   data_col74[19] <= data_col74[18];
   data_col74[20] <= data_col74[19];
   data_col74[21] <= data_col74[20];
   data_col74[22] <= data_col74[21];
   data_col74[23] <= data_col74[22];
   data_col74[24] <= data_col74[23];
   data_col74[25] <= data_col74[24];
   data_col74[26] <= data_col74[25];
   data_col74[27] <= data_col74[26];
   data_col74[28] <= data_col74[27];
   data_col74[29] <= data_col74[28];
   data_col74[30] <= data_col74[29];
   data_col74[31] <= data_col74[30];
   data_col74[32] <= data_col74[31];
   data_col74[33] <= data_col74[32];
   data_col74[34] <= data_col74[33];
   data_col74[35] <= data_col74[34];
   data_col74[36] <= data_col74[35];
   data_col74[37] <= data_col74[36];
   data_col74[38] <= data_col74[37];
   data_col74[39] <= data_col74[38];
   data_col74[40] <= data_col74[39];
   data_col74[41] <= data_col74[40];
   data_col74[42] <= data_col74[41];
   data_col74[43] <= data_col74[42];
   data_col74[44] <= data_col74[43];
   data_col74[45] <= data_col74[44];
   data_col74[46] <= data_col74[45];
   data_col74[47] <= data_col74[46];
   data_col74[48] <= data_col74[47];
   data_col74[49] <= data_col74[48];
   data_col74[50] <= data_col74[49];
   data_col74[51] <= data_col74[50];
   data_col74[52] <= data_col74[51];
   data_col74[53] <= data_col74[52];
   data_col74[54] <= data_col74[53];
   data_col74[55] <= data_col74[54];
   data_col74[56] <= data_col74[55];
   data_col74[57] <= data_col74[56];
   data_col74[58] <= data_col74[57];
   data_col74[59] <= data_col74[58];
   data_col74[60] <= data_col74[59];
   data_col74[61] <= data_col74[60];
   data_col74[62] <= data_col74[61];
   data_col74[63] <= data_col74[62];
   data_col74[64] <= data_col74[63];
   data_col74[65] <= data_col74[64];
   data_col74[66] <= data_col74[65];
   data_col74[67] <= data_col74[66];
   data_col74[68] <= data_col74[67];
   data_col74[69] <= data_col74[68];
   data_col74[70] <= data_col74[69];
   data_col74[71] <= data_col74[70];
   data_col74[72] <= data_col74[71];
   data_col74[73] <= data_col74[72];
   data_col74[74] <= data_col74[73];

   data_col75[1] <= data[25];
   data_col75[2] <= data_col75[1];
   data_col75[3] <= data_col75[2];
   data_col75[4] <= data_col75[3];
   data_col75[5] <= data_col75[4];
   data_col75[6] <= data_col75[5];
   data_col75[7] <= data_col75[6];
   data_col75[8] <= data_col75[7];
   data_col75[9] <= data_col75[8];
   data_col75[10] <= data_col75[9];
   data_col75[11] <= data_col75[10];
   data_col75[12] <= data_col75[11];
   data_col75[13] <= data_col75[12];
   data_col75[14] <= data_col75[13];
   data_col75[15] <= data_col75[14];
   data_col75[16] <= data_col75[15];
   data_col75[17] <= data_col75[16];
   data_col75[18] <= data_col75[17];
   data_col75[19] <= data_col75[18];
   data_col75[20] <= data_col75[19];
   data_col75[21] <= data_col75[20];
   data_col75[22] <= data_col75[21];
   data_col75[23] <= data_col75[22];
   data_col75[24] <= data_col75[23];
   data_col75[25] <= data_col75[24];
   data_col75[26] <= data_col75[25];
   data_col75[27] <= data_col75[26];
   data_col75[28] <= data_col75[27];
   data_col75[29] <= data_col75[28];
   data_col75[30] <= data_col75[29];
   data_col75[31] <= data_col75[30];
   data_col75[32] <= data_col75[31];
   data_col75[33] <= data_col75[32];
   data_col75[34] <= data_col75[33];
   data_col75[35] <= data_col75[34];
   data_col75[36] <= data_col75[35];
   data_col75[37] <= data_col75[36];
   data_col75[38] <= data_col75[37];
   data_col75[39] <= data_col75[38];
   data_col75[40] <= data_col75[39];
   data_col75[41] <= data_col75[40];
   data_col75[42] <= data_col75[41];
   data_col75[43] <= data_col75[42];
   data_col75[44] <= data_col75[43];
   data_col75[45] <= data_col75[44];
   data_col75[46] <= data_col75[45];
   data_col75[47] <= data_col75[46];
   data_col75[48] <= data_col75[47];
   data_col75[49] <= data_col75[48];
   data_col75[50] <= data_col75[49];
   data_col75[51] <= data_col75[50];
   data_col75[52] <= data_col75[51];
   data_col75[53] <= data_col75[52];
   data_col75[54] <= data_col75[53];
   data_col75[55] <= data_col75[54];
   data_col75[56] <= data_col75[55];
   data_col75[57] <= data_col75[56];
   data_col75[58] <= data_col75[57];
   data_col75[59] <= data_col75[58];
   data_col75[60] <= data_col75[59];
   data_col75[61] <= data_col75[60];
   data_col75[62] <= data_col75[61];
   data_col75[63] <= data_col75[62];
   data_col75[64] <= data_col75[63];
   data_col75[65] <= data_col75[64];
   data_col75[66] <= data_col75[65];
   data_col75[67] <= data_col75[66];
   data_col75[68] <= data_col75[67];
   data_col75[69] <= data_col75[68];
   data_col75[70] <= data_col75[69];
   data_col75[71] <= data_col75[70];
   data_col75[72] <= data_col75[71];
   data_col75[73] <= data_col75[72];
   data_col75[74] <= data_col75[73];
   data_col75[75] <= data_col75[74];

   data_col76[1] <= data[24];
   data_col76[2] <= data_col76[1];
   data_col76[3] <= data_col76[2];
   data_col76[4] <= data_col76[3];
   data_col76[5] <= data_col76[4];
   data_col76[6] <= data_col76[5];
   data_col76[7] <= data_col76[6];
   data_col76[8] <= data_col76[7];
   data_col76[9] <= data_col76[8];
   data_col76[10] <= data_col76[9];
   data_col76[11] <= data_col76[10];
   data_col76[12] <= data_col76[11];
   data_col76[13] <= data_col76[12];
   data_col76[14] <= data_col76[13];
   data_col76[15] <= data_col76[14];
   data_col76[16] <= data_col76[15];
   data_col76[17] <= data_col76[16];
   data_col76[18] <= data_col76[17];
   data_col76[19] <= data_col76[18];
   data_col76[20] <= data_col76[19];
   data_col76[21] <= data_col76[20];
   data_col76[22] <= data_col76[21];
   data_col76[23] <= data_col76[22];
   data_col76[24] <= data_col76[23];
   data_col76[25] <= data_col76[24];
   data_col76[26] <= data_col76[25];
   data_col76[27] <= data_col76[26];
   data_col76[28] <= data_col76[27];
   data_col76[29] <= data_col76[28];
   data_col76[30] <= data_col76[29];
   data_col76[31] <= data_col76[30];
   data_col76[32] <= data_col76[31];
   data_col76[33] <= data_col76[32];
   data_col76[34] <= data_col76[33];
   data_col76[35] <= data_col76[34];
   data_col76[36] <= data_col76[35];
   data_col76[37] <= data_col76[36];
   data_col76[38] <= data_col76[37];
   data_col76[39] <= data_col76[38];
   data_col76[40] <= data_col76[39];
   data_col76[41] <= data_col76[40];
   data_col76[42] <= data_col76[41];
   data_col76[43] <= data_col76[42];
   data_col76[44] <= data_col76[43];
   data_col76[45] <= data_col76[44];
   data_col76[46] <= data_col76[45];
   data_col76[47] <= data_col76[46];
   data_col76[48] <= data_col76[47];
   data_col76[49] <= data_col76[48];
   data_col76[50] <= data_col76[49];
   data_col76[51] <= data_col76[50];
   data_col76[52] <= data_col76[51];
   data_col76[53] <= data_col76[52];
   data_col76[54] <= data_col76[53];
   data_col76[55] <= data_col76[54];
   data_col76[56] <= data_col76[55];
   data_col76[57] <= data_col76[56];
   data_col76[58] <= data_col76[57];
   data_col76[59] <= data_col76[58];
   data_col76[60] <= data_col76[59];
   data_col76[61] <= data_col76[60];
   data_col76[62] <= data_col76[61];
   data_col76[63] <= data_col76[62];
   data_col76[64] <= data_col76[63];
   data_col76[65] <= data_col76[64];
   data_col76[66] <= data_col76[65];
   data_col76[67] <= data_col76[66];
   data_col76[68] <= data_col76[67];
   data_col76[69] <= data_col76[68];
   data_col76[70] <= data_col76[69];
   data_col76[71] <= data_col76[70];
   data_col76[72] <= data_col76[71];
   data_col76[73] <= data_col76[72];
   data_col76[74] <= data_col76[73];
   data_col76[75] <= data_col76[74];
   data_col76[76] <= data_col76[75];

   data_col77[1] <= data[23];
   data_col77[2] <= data_col77[1];
   data_col77[3] <= data_col77[2];
   data_col77[4] <= data_col77[3];
   data_col77[5] <= data_col77[4];
   data_col77[6] <= data_col77[5];
   data_col77[7] <= data_col77[6];
   data_col77[8] <= data_col77[7];
   data_col77[9] <= data_col77[8];
   data_col77[10] <= data_col77[9];
   data_col77[11] <= data_col77[10];
   data_col77[12] <= data_col77[11];
   data_col77[13] <= data_col77[12];
   data_col77[14] <= data_col77[13];
   data_col77[15] <= data_col77[14];
   data_col77[16] <= data_col77[15];
   data_col77[17] <= data_col77[16];
   data_col77[18] <= data_col77[17];
   data_col77[19] <= data_col77[18];
   data_col77[20] <= data_col77[19];
   data_col77[21] <= data_col77[20];
   data_col77[22] <= data_col77[21];
   data_col77[23] <= data_col77[22];
   data_col77[24] <= data_col77[23];
   data_col77[25] <= data_col77[24];
   data_col77[26] <= data_col77[25];
   data_col77[27] <= data_col77[26];
   data_col77[28] <= data_col77[27];
   data_col77[29] <= data_col77[28];
   data_col77[30] <= data_col77[29];
   data_col77[31] <= data_col77[30];
   data_col77[32] <= data_col77[31];
   data_col77[33] <= data_col77[32];
   data_col77[34] <= data_col77[33];
   data_col77[35] <= data_col77[34];
   data_col77[36] <= data_col77[35];
   data_col77[37] <= data_col77[36];
   data_col77[38] <= data_col77[37];
   data_col77[39] <= data_col77[38];
   data_col77[40] <= data_col77[39];
   data_col77[41] <= data_col77[40];
   data_col77[42] <= data_col77[41];
   data_col77[43] <= data_col77[42];
   data_col77[44] <= data_col77[43];
   data_col77[45] <= data_col77[44];
   data_col77[46] <= data_col77[45];
   data_col77[47] <= data_col77[46];
   data_col77[48] <= data_col77[47];
   data_col77[49] <= data_col77[48];
   data_col77[50] <= data_col77[49];
   data_col77[51] <= data_col77[50];
   data_col77[52] <= data_col77[51];
   data_col77[53] <= data_col77[52];
   data_col77[54] <= data_col77[53];
   data_col77[55] <= data_col77[54];
   data_col77[56] <= data_col77[55];
   data_col77[57] <= data_col77[56];
   data_col77[58] <= data_col77[57];
   data_col77[59] <= data_col77[58];
   data_col77[60] <= data_col77[59];
   data_col77[61] <= data_col77[60];
   data_col77[62] <= data_col77[61];
   data_col77[63] <= data_col77[62];
   data_col77[64] <= data_col77[63];
   data_col77[65] <= data_col77[64];
   data_col77[66] <= data_col77[65];
   data_col77[67] <= data_col77[66];
   data_col77[68] <= data_col77[67];
   data_col77[69] <= data_col77[68];
   data_col77[70] <= data_col77[69];
   data_col77[71] <= data_col77[70];
   data_col77[72] <= data_col77[71];
   data_col77[73] <= data_col77[72];
   data_col77[74] <= data_col77[73];
   data_col77[75] <= data_col77[74];
   data_col77[76] <= data_col77[75];
   data_col77[77] <= data_col77[76];

   data_col78[1] <= data[22];
   data_col78[2] <= data_col78[1];
   data_col78[3] <= data_col78[2];
   data_col78[4] <= data_col78[3];
   data_col78[5] <= data_col78[4];
   data_col78[6] <= data_col78[5];
   data_col78[7] <= data_col78[6];
   data_col78[8] <= data_col78[7];
   data_col78[9] <= data_col78[8];
   data_col78[10] <= data_col78[9];
   data_col78[11] <= data_col78[10];
   data_col78[12] <= data_col78[11];
   data_col78[13] <= data_col78[12];
   data_col78[14] <= data_col78[13];
   data_col78[15] <= data_col78[14];
   data_col78[16] <= data_col78[15];
   data_col78[17] <= data_col78[16];
   data_col78[18] <= data_col78[17];
   data_col78[19] <= data_col78[18];
   data_col78[20] <= data_col78[19];
   data_col78[21] <= data_col78[20];
   data_col78[22] <= data_col78[21];
   data_col78[23] <= data_col78[22];
   data_col78[24] <= data_col78[23];
   data_col78[25] <= data_col78[24];
   data_col78[26] <= data_col78[25];
   data_col78[27] <= data_col78[26];
   data_col78[28] <= data_col78[27];
   data_col78[29] <= data_col78[28];
   data_col78[30] <= data_col78[29];
   data_col78[31] <= data_col78[30];
   data_col78[32] <= data_col78[31];
   data_col78[33] <= data_col78[32];
   data_col78[34] <= data_col78[33];
   data_col78[35] <= data_col78[34];
   data_col78[36] <= data_col78[35];
   data_col78[37] <= data_col78[36];
   data_col78[38] <= data_col78[37];
   data_col78[39] <= data_col78[38];
   data_col78[40] <= data_col78[39];
   data_col78[41] <= data_col78[40];
   data_col78[42] <= data_col78[41];
   data_col78[43] <= data_col78[42];
   data_col78[44] <= data_col78[43];
   data_col78[45] <= data_col78[44];
   data_col78[46] <= data_col78[45];
   data_col78[47] <= data_col78[46];
   data_col78[48] <= data_col78[47];
   data_col78[49] <= data_col78[48];
   data_col78[50] <= data_col78[49];
   data_col78[51] <= data_col78[50];
   data_col78[52] <= data_col78[51];
   data_col78[53] <= data_col78[52];
   data_col78[54] <= data_col78[53];
   data_col78[55] <= data_col78[54];
   data_col78[56] <= data_col78[55];
   data_col78[57] <= data_col78[56];
   data_col78[58] <= data_col78[57];
   data_col78[59] <= data_col78[58];
   data_col78[60] <= data_col78[59];
   data_col78[61] <= data_col78[60];
   data_col78[62] <= data_col78[61];
   data_col78[63] <= data_col78[62];
   data_col78[64] <= data_col78[63];
   data_col78[65] <= data_col78[64];
   data_col78[66] <= data_col78[65];
   data_col78[67] <= data_col78[66];
   data_col78[68] <= data_col78[67];
   data_col78[69] <= data_col78[68];
   data_col78[70] <= data_col78[69];
   data_col78[71] <= data_col78[70];
   data_col78[72] <= data_col78[71];
   data_col78[73] <= data_col78[72];
   data_col78[74] <= data_col78[73];
   data_col78[75] <= data_col78[74];
   data_col78[76] <= data_col78[75];
   data_col78[77] <= data_col78[76];
   data_col78[78] <= data_col78[77];

   data_col79[1] <= data[21];
   data_col79[2] <= data_col79[1];
   data_col79[3] <= data_col79[2];
   data_col79[4] <= data_col79[3];
   data_col79[5] <= data_col79[4];
   data_col79[6] <= data_col79[5];
   data_col79[7] <= data_col79[6];
   data_col79[8] <= data_col79[7];
   data_col79[9] <= data_col79[8];
   data_col79[10] <= data_col79[9];
   data_col79[11] <= data_col79[10];
   data_col79[12] <= data_col79[11];
   data_col79[13] <= data_col79[12];
   data_col79[14] <= data_col79[13];
   data_col79[15] <= data_col79[14];
   data_col79[16] <= data_col79[15];
   data_col79[17] <= data_col79[16];
   data_col79[18] <= data_col79[17];
   data_col79[19] <= data_col79[18];
   data_col79[20] <= data_col79[19];
   data_col79[21] <= data_col79[20];
   data_col79[22] <= data_col79[21];
   data_col79[23] <= data_col79[22];
   data_col79[24] <= data_col79[23];
   data_col79[25] <= data_col79[24];
   data_col79[26] <= data_col79[25];
   data_col79[27] <= data_col79[26];
   data_col79[28] <= data_col79[27];
   data_col79[29] <= data_col79[28];
   data_col79[30] <= data_col79[29];
   data_col79[31] <= data_col79[30];
   data_col79[32] <= data_col79[31];
   data_col79[33] <= data_col79[32];
   data_col79[34] <= data_col79[33];
   data_col79[35] <= data_col79[34];
   data_col79[36] <= data_col79[35];
   data_col79[37] <= data_col79[36];
   data_col79[38] <= data_col79[37];
   data_col79[39] <= data_col79[38];
   data_col79[40] <= data_col79[39];
   data_col79[41] <= data_col79[40];
   data_col79[42] <= data_col79[41];
   data_col79[43] <= data_col79[42];
   data_col79[44] <= data_col79[43];
   data_col79[45] <= data_col79[44];
   data_col79[46] <= data_col79[45];
   data_col79[47] <= data_col79[46];
   data_col79[48] <= data_col79[47];
   data_col79[49] <= data_col79[48];
   data_col79[50] <= data_col79[49];
   data_col79[51] <= data_col79[50];
   data_col79[52] <= data_col79[51];
   data_col79[53] <= data_col79[52];
   data_col79[54] <= data_col79[53];
   data_col79[55] <= data_col79[54];
   data_col79[56] <= data_col79[55];
   data_col79[57] <= data_col79[56];
   data_col79[58] <= data_col79[57];
   data_col79[59] <= data_col79[58];
   data_col79[60] <= data_col79[59];
   data_col79[61] <= data_col79[60];
   data_col79[62] <= data_col79[61];
   data_col79[63] <= data_col79[62];
   data_col79[64] <= data_col79[63];
   data_col79[65] <= data_col79[64];
   data_col79[66] <= data_col79[65];
   data_col79[67] <= data_col79[66];
   data_col79[68] <= data_col79[67];
   data_col79[69] <= data_col79[68];
   data_col79[70] <= data_col79[69];
   data_col79[71] <= data_col79[70];
   data_col79[72] <= data_col79[71];
   data_col79[73] <= data_col79[72];
   data_col79[74] <= data_col79[73];
   data_col79[75] <= data_col79[74];
   data_col79[76] <= data_col79[75];
   data_col79[77] <= data_col79[76];
   data_col79[78] <= data_col79[77];
   data_col79[79] <= data_col79[78];

   data_col80[1] <= data[20];
   data_col80[2] <= data_col80[1];
   data_col80[3] <= data_col80[2];
   data_col80[4] <= data_col80[3];
   data_col80[5] <= data_col80[4];
   data_col80[6] <= data_col80[5];
   data_col80[7] <= data_col80[6];
   data_col80[8] <= data_col80[7];
   data_col80[9] <= data_col80[8];
   data_col80[10] <= data_col80[9];
   data_col80[11] <= data_col80[10];
   data_col80[12] <= data_col80[11];
   data_col80[13] <= data_col80[12];
   data_col80[14] <= data_col80[13];
   data_col80[15] <= data_col80[14];
   data_col80[16] <= data_col80[15];
   data_col80[17] <= data_col80[16];
   data_col80[18] <= data_col80[17];
   data_col80[19] <= data_col80[18];
   data_col80[20] <= data_col80[19];
   data_col80[21] <= data_col80[20];
   data_col80[22] <= data_col80[21];
   data_col80[23] <= data_col80[22];
   data_col80[24] <= data_col80[23];
   data_col80[25] <= data_col80[24];
   data_col80[26] <= data_col80[25];
   data_col80[27] <= data_col80[26];
   data_col80[28] <= data_col80[27];
   data_col80[29] <= data_col80[28];
   data_col80[30] <= data_col80[29];
   data_col80[31] <= data_col80[30];
   data_col80[32] <= data_col80[31];
   data_col80[33] <= data_col80[32];
   data_col80[34] <= data_col80[33];
   data_col80[35] <= data_col80[34];
   data_col80[36] <= data_col80[35];
   data_col80[37] <= data_col80[36];
   data_col80[38] <= data_col80[37];
   data_col80[39] <= data_col80[38];
   data_col80[40] <= data_col80[39];
   data_col80[41] <= data_col80[40];
   data_col80[42] <= data_col80[41];
   data_col80[43] <= data_col80[42];
   data_col80[44] <= data_col80[43];
   data_col80[45] <= data_col80[44];
   data_col80[46] <= data_col80[45];
   data_col80[47] <= data_col80[46];
   data_col80[48] <= data_col80[47];
   data_col80[49] <= data_col80[48];
   data_col80[50] <= data_col80[49];
   data_col80[51] <= data_col80[50];
   data_col80[52] <= data_col80[51];
   data_col80[53] <= data_col80[52];
   data_col80[54] <= data_col80[53];
   data_col80[55] <= data_col80[54];
   data_col80[56] <= data_col80[55];
   data_col80[57] <= data_col80[56];
   data_col80[58] <= data_col80[57];
   data_col80[59] <= data_col80[58];
   data_col80[60] <= data_col80[59];
   data_col80[61] <= data_col80[60];
   data_col80[62] <= data_col80[61];
   data_col80[63] <= data_col80[62];
   data_col80[64] <= data_col80[63];
   data_col80[65] <= data_col80[64];
   data_col80[66] <= data_col80[65];
   data_col80[67] <= data_col80[66];
   data_col80[68] <= data_col80[67];
   data_col80[69] <= data_col80[68];
   data_col80[70] <= data_col80[69];
   data_col80[71] <= data_col80[70];
   data_col80[72] <= data_col80[71];
   data_col80[73] <= data_col80[72];
   data_col80[74] <= data_col80[73];
   data_col80[75] <= data_col80[74];
   data_col80[76] <= data_col80[75];
   data_col80[77] <= data_col80[76];
   data_col80[78] <= data_col80[77];
   data_col80[79] <= data_col80[78];
   data_col80[80] <= data_col80[79];

   data_col81[1] <= data[19];
   data_col81[2] <= data_col81[1];
   data_col81[3] <= data_col81[2];
   data_col81[4] <= data_col81[3];
   data_col81[5] <= data_col81[4];
   data_col81[6] <= data_col81[5];
   data_col81[7] <= data_col81[6];
   data_col81[8] <= data_col81[7];
   data_col81[9] <= data_col81[8];
   data_col81[10] <= data_col81[9];
   data_col81[11] <= data_col81[10];
   data_col81[12] <= data_col81[11];
   data_col81[13] <= data_col81[12];
   data_col81[14] <= data_col81[13];
   data_col81[15] <= data_col81[14];
   data_col81[16] <= data_col81[15];
   data_col81[17] <= data_col81[16];
   data_col81[18] <= data_col81[17];
   data_col81[19] <= data_col81[18];
   data_col81[20] <= data_col81[19];
   data_col81[21] <= data_col81[20];
   data_col81[22] <= data_col81[21];
   data_col81[23] <= data_col81[22];
   data_col81[24] <= data_col81[23];
   data_col81[25] <= data_col81[24];
   data_col81[26] <= data_col81[25];
   data_col81[27] <= data_col81[26];
   data_col81[28] <= data_col81[27];
   data_col81[29] <= data_col81[28];
   data_col81[30] <= data_col81[29];
   data_col81[31] <= data_col81[30];
   data_col81[32] <= data_col81[31];
   data_col81[33] <= data_col81[32];
   data_col81[34] <= data_col81[33];
   data_col81[35] <= data_col81[34];
   data_col81[36] <= data_col81[35];
   data_col81[37] <= data_col81[36];
   data_col81[38] <= data_col81[37];
   data_col81[39] <= data_col81[38];
   data_col81[40] <= data_col81[39];
   data_col81[41] <= data_col81[40];
   data_col81[42] <= data_col81[41];
   data_col81[43] <= data_col81[42];
   data_col81[44] <= data_col81[43];
   data_col81[45] <= data_col81[44];
   data_col81[46] <= data_col81[45];
   data_col81[47] <= data_col81[46];
   data_col81[48] <= data_col81[47];
   data_col81[49] <= data_col81[48];
   data_col81[50] <= data_col81[49];
   data_col81[51] <= data_col81[50];
   data_col81[52] <= data_col81[51];
   data_col81[53] <= data_col81[52];
   data_col81[54] <= data_col81[53];
   data_col81[55] <= data_col81[54];
   data_col81[56] <= data_col81[55];
   data_col81[57] <= data_col81[56];
   data_col81[58] <= data_col81[57];
   data_col81[59] <= data_col81[58];
   data_col81[60] <= data_col81[59];
   data_col81[61] <= data_col81[60];
   data_col81[62] <= data_col81[61];
   data_col81[63] <= data_col81[62];
   data_col81[64] <= data_col81[63];
   data_col81[65] <= data_col81[64];
   data_col81[66] <= data_col81[65];
   data_col81[67] <= data_col81[66];
   data_col81[68] <= data_col81[67];
   data_col81[69] <= data_col81[68];
   data_col81[70] <= data_col81[69];
   data_col81[71] <= data_col81[70];
   data_col81[72] <= data_col81[71];
   data_col81[73] <= data_col81[72];
   data_col81[74] <= data_col81[73];
   data_col81[75] <= data_col81[74];
   data_col81[76] <= data_col81[75];
   data_col81[77] <= data_col81[76];
   data_col81[78] <= data_col81[77];
   data_col81[79] <= data_col81[78];
   data_col81[80] <= data_col81[79];
   data_col81[81] <= data_col81[80];

   data_col82[1] <= data[18];
   data_col82[2] <= data_col82[1];
   data_col82[3] <= data_col82[2];
   data_col82[4] <= data_col82[3];
   data_col82[5] <= data_col82[4];
   data_col82[6] <= data_col82[5];
   data_col82[7] <= data_col82[6];
   data_col82[8] <= data_col82[7];
   data_col82[9] <= data_col82[8];
   data_col82[10] <= data_col82[9];
   data_col82[11] <= data_col82[10];
   data_col82[12] <= data_col82[11];
   data_col82[13] <= data_col82[12];
   data_col82[14] <= data_col82[13];
   data_col82[15] <= data_col82[14];
   data_col82[16] <= data_col82[15];
   data_col82[17] <= data_col82[16];
   data_col82[18] <= data_col82[17];
   data_col82[19] <= data_col82[18];
   data_col82[20] <= data_col82[19];
   data_col82[21] <= data_col82[20];
   data_col82[22] <= data_col82[21];
   data_col82[23] <= data_col82[22];
   data_col82[24] <= data_col82[23];
   data_col82[25] <= data_col82[24];
   data_col82[26] <= data_col82[25];
   data_col82[27] <= data_col82[26];
   data_col82[28] <= data_col82[27];
   data_col82[29] <= data_col82[28];
   data_col82[30] <= data_col82[29];
   data_col82[31] <= data_col82[30];
   data_col82[32] <= data_col82[31];
   data_col82[33] <= data_col82[32];
   data_col82[34] <= data_col82[33];
   data_col82[35] <= data_col82[34];
   data_col82[36] <= data_col82[35];
   data_col82[37] <= data_col82[36];
   data_col82[38] <= data_col82[37];
   data_col82[39] <= data_col82[38];
   data_col82[40] <= data_col82[39];
   data_col82[41] <= data_col82[40];
   data_col82[42] <= data_col82[41];
   data_col82[43] <= data_col82[42];
   data_col82[44] <= data_col82[43];
   data_col82[45] <= data_col82[44];
   data_col82[46] <= data_col82[45];
   data_col82[47] <= data_col82[46];
   data_col82[48] <= data_col82[47];
   data_col82[49] <= data_col82[48];
   data_col82[50] <= data_col82[49];
   data_col82[51] <= data_col82[50];
   data_col82[52] <= data_col82[51];
   data_col82[53] <= data_col82[52];
   data_col82[54] <= data_col82[53];
   data_col82[55] <= data_col82[54];
   data_col82[56] <= data_col82[55];
   data_col82[57] <= data_col82[56];
   data_col82[58] <= data_col82[57];
   data_col82[59] <= data_col82[58];
   data_col82[60] <= data_col82[59];
   data_col82[61] <= data_col82[60];
   data_col82[62] <= data_col82[61];
   data_col82[63] <= data_col82[62];
   data_col82[64] <= data_col82[63];
   data_col82[65] <= data_col82[64];
   data_col82[66] <= data_col82[65];
   data_col82[67] <= data_col82[66];
   data_col82[68] <= data_col82[67];
   data_col82[69] <= data_col82[68];
   data_col82[70] <= data_col82[69];
   data_col82[71] <= data_col82[70];
   data_col82[72] <= data_col82[71];
   data_col82[73] <= data_col82[72];
   data_col82[74] <= data_col82[73];
   data_col82[75] <= data_col82[74];
   data_col82[76] <= data_col82[75];
   data_col82[77] <= data_col82[76];
   data_col82[78] <= data_col82[77];
   data_col82[79] <= data_col82[78];
   data_col82[80] <= data_col82[79];
   data_col82[81] <= data_col82[80];
   data_col82[82] <= data_col82[81];

   data_col83[1] <= data[17];
   data_col83[2] <= data_col83[1];
   data_col83[3] <= data_col83[2];
   data_col83[4] <= data_col83[3];
   data_col83[5] <= data_col83[4];
   data_col83[6] <= data_col83[5];
   data_col83[7] <= data_col83[6];
   data_col83[8] <= data_col83[7];
   data_col83[9] <= data_col83[8];
   data_col83[10] <= data_col83[9];
   data_col83[11] <= data_col83[10];
   data_col83[12] <= data_col83[11];
   data_col83[13] <= data_col83[12];
   data_col83[14] <= data_col83[13];
   data_col83[15] <= data_col83[14];
   data_col83[16] <= data_col83[15];
   data_col83[17] <= data_col83[16];
   data_col83[18] <= data_col83[17];
   data_col83[19] <= data_col83[18];
   data_col83[20] <= data_col83[19];
   data_col83[21] <= data_col83[20];
   data_col83[22] <= data_col83[21];
   data_col83[23] <= data_col83[22];
   data_col83[24] <= data_col83[23];
   data_col83[25] <= data_col83[24];
   data_col83[26] <= data_col83[25];
   data_col83[27] <= data_col83[26];
   data_col83[28] <= data_col83[27];
   data_col83[29] <= data_col83[28];
   data_col83[30] <= data_col83[29];
   data_col83[31] <= data_col83[30];
   data_col83[32] <= data_col83[31];
   data_col83[33] <= data_col83[32];
   data_col83[34] <= data_col83[33];
   data_col83[35] <= data_col83[34];
   data_col83[36] <= data_col83[35];
   data_col83[37] <= data_col83[36];
   data_col83[38] <= data_col83[37];
   data_col83[39] <= data_col83[38];
   data_col83[40] <= data_col83[39];
   data_col83[41] <= data_col83[40];
   data_col83[42] <= data_col83[41];
   data_col83[43] <= data_col83[42];
   data_col83[44] <= data_col83[43];
   data_col83[45] <= data_col83[44];
   data_col83[46] <= data_col83[45];
   data_col83[47] <= data_col83[46];
   data_col83[48] <= data_col83[47];
   data_col83[49] <= data_col83[48];
   data_col83[50] <= data_col83[49];
   data_col83[51] <= data_col83[50];
   data_col83[52] <= data_col83[51];
   data_col83[53] <= data_col83[52];
   data_col83[54] <= data_col83[53];
   data_col83[55] <= data_col83[54];
   data_col83[56] <= data_col83[55];
   data_col83[57] <= data_col83[56];
   data_col83[58] <= data_col83[57];
   data_col83[59] <= data_col83[58];
   data_col83[60] <= data_col83[59];
   data_col83[61] <= data_col83[60];
   data_col83[62] <= data_col83[61];
   data_col83[63] <= data_col83[62];
   data_col83[64] <= data_col83[63];
   data_col83[65] <= data_col83[64];
   data_col83[66] <= data_col83[65];
   data_col83[67] <= data_col83[66];
   data_col83[68] <= data_col83[67];
   data_col83[69] <= data_col83[68];
   data_col83[70] <= data_col83[69];
   data_col83[71] <= data_col83[70];
   data_col83[72] <= data_col83[71];
   data_col83[73] <= data_col83[72];
   data_col83[74] <= data_col83[73];
   data_col83[75] <= data_col83[74];
   data_col83[76] <= data_col83[75];
   data_col83[77] <= data_col83[76];
   data_col83[78] <= data_col83[77];
   data_col83[79] <= data_col83[78];
   data_col83[80] <= data_col83[79];
   data_col83[81] <= data_col83[80];
   data_col83[82] <= data_col83[81];
   data_col83[83] <= data_col83[82];

   data_col84[1] <= data[16];
   data_col84[2] <= data_col84[1];
   data_col84[3] <= data_col84[2];
   data_col84[4] <= data_col84[3];
   data_col84[5] <= data_col84[4];
   data_col84[6] <= data_col84[5];
   data_col84[7] <= data_col84[6];
   data_col84[8] <= data_col84[7];
   data_col84[9] <= data_col84[8];
   data_col84[10] <= data_col84[9];
   data_col84[11] <= data_col84[10];
   data_col84[12] <= data_col84[11];
   data_col84[13] <= data_col84[12];
   data_col84[14] <= data_col84[13];
   data_col84[15] <= data_col84[14];
   data_col84[16] <= data_col84[15];
   data_col84[17] <= data_col84[16];
   data_col84[18] <= data_col84[17];
   data_col84[19] <= data_col84[18];
   data_col84[20] <= data_col84[19];
   data_col84[21] <= data_col84[20];
   data_col84[22] <= data_col84[21];
   data_col84[23] <= data_col84[22];
   data_col84[24] <= data_col84[23];
   data_col84[25] <= data_col84[24];
   data_col84[26] <= data_col84[25];
   data_col84[27] <= data_col84[26];
   data_col84[28] <= data_col84[27];
   data_col84[29] <= data_col84[28];
   data_col84[30] <= data_col84[29];
   data_col84[31] <= data_col84[30];
   data_col84[32] <= data_col84[31];
   data_col84[33] <= data_col84[32];
   data_col84[34] <= data_col84[33];
   data_col84[35] <= data_col84[34];
   data_col84[36] <= data_col84[35];
   data_col84[37] <= data_col84[36];
   data_col84[38] <= data_col84[37];
   data_col84[39] <= data_col84[38];
   data_col84[40] <= data_col84[39];
   data_col84[41] <= data_col84[40];
   data_col84[42] <= data_col84[41];
   data_col84[43] <= data_col84[42];
   data_col84[44] <= data_col84[43];
   data_col84[45] <= data_col84[44];
   data_col84[46] <= data_col84[45];
   data_col84[47] <= data_col84[46];
   data_col84[48] <= data_col84[47];
   data_col84[49] <= data_col84[48];
   data_col84[50] <= data_col84[49];
   data_col84[51] <= data_col84[50];
   data_col84[52] <= data_col84[51];
   data_col84[53] <= data_col84[52];
   data_col84[54] <= data_col84[53];
   data_col84[55] <= data_col84[54];
   data_col84[56] <= data_col84[55];
   data_col84[57] <= data_col84[56];
   data_col84[58] <= data_col84[57];
   data_col84[59] <= data_col84[58];
   data_col84[60] <= data_col84[59];
   data_col84[61] <= data_col84[60];
   data_col84[62] <= data_col84[61];
   data_col84[63] <= data_col84[62];
   data_col84[64] <= data_col84[63];
   data_col84[65] <= data_col84[64];
   data_col84[66] <= data_col84[65];
   data_col84[67] <= data_col84[66];
   data_col84[68] <= data_col84[67];
   data_col84[69] <= data_col84[68];
   data_col84[70] <= data_col84[69];
   data_col84[71] <= data_col84[70];
   data_col84[72] <= data_col84[71];
   data_col84[73] <= data_col84[72];
   data_col84[74] <= data_col84[73];
   data_col84[75] <= data_col84[74];
   data_col84[76] <= data_col84[75];
   data_col84[77] <= data_col84[76];
   data_col84[78] <= data_col84[77];
   data_col84[79] <= data_col84[78];
   data_col84[80] <= data_col84[79];
   data_col84[81] <= data_col84[80];
   data_col84[82] <= data_col84[81];
   data_col84[83] <= data_col84[82];
   data_col84[84] <= data_col84[83];

   data_col85[1] <= data[15];
   data_col85[2] <= data_col85[1];
   data_col85[3] <= data_col85[2];
   data_col85[4] <= data_col85[3];
   data_col85[5] <= data_col85[4];
   data_col85[6] <= data_col85[5];
   data_col85[7] <= data_col85[6];
   data_col85[8] <= data_col85[7];
   data_col85[9] <= data_col85[8];
   data_col85[10] <= data_col85[9];
   data_col85[11] <= data_col85[10];
   data_col85[12] <= data_col85[11];
   data_col85[13] <= data_col85[12];
   data_col85[14] <= data_col85[13];
   data_col85[15] <= data_col85[14];
   data_col85[16] <= data_col85[15];
   data_col85[17] <= data_col85[16];
   data_col85[18] <= data_col85[17];
   data_col85[19] <= data_col85[18];
   data_col85[20] <= data_col85[19];
   data_col85[21] <= data_col85[20];
   data_col85[22] <= data_col85[21];
   data_col85[23] <= data_col85[22];
   data_col85[24] <= data_col85[23];
   data_col85[25] <= data_col85[24];
   data_col85[26] <= data_col85[25];
   data_col85[27] <= data_col85[26];
   data_col85[28] <= data_col85[27];
   data_col85[29] <= data_col85[28];
   data_col85[30] <= data_col85[29];
   data_col85[31] <= data_col85[30];
   data_col85[32] <= data_col85[31];
   data_col85[33] <= data_col85[32];
   data_col85[34] <= data_col85[33];
   data_col85[35] <= data_col85[34];
   data_col85[36] <= data_col85[35];
   data_col85[37] <= data_col85[36];
   data_col85[38] <= data_col85[37];
   data_col85[39] <= data_col85[38];
   data_col85[40] <= data_col85[39];
   data_col85[41] <= data_col85[40];
   data_col85[42] <= data_col85[41];
   data_col85[43] <= data_col85[42];
   data_col85[44] <= data_col85[43];
   data_col85[45] <= data_col85[44];
   data_col85[46] <= data_col85[45];
   data_col85[47] <= data_col85[46];
   data_col85[48] <= data_col85[47];
   data_col85[49] <= data_col85[48];
   data_col85[50] <= data_col85[49];
   data_col85[51] <= data_col85[50];
   data_col85[52] <= data_col85[51];
   data_col85[53] <= data_col85[52];
   data_col85[54] <= data_col85[53];
   data_col85[55] <= data_col85[54];
   data_col85[56] <= data_col85[55];
   data_col85[57] <= data_col85[56];
   data_col85[58] <= data_col85[57];
   data_col85[59] <= data_col85[58];
   data_col85[60] <= data_col85[59];
   data_col85[61] <= data_col85[60];
   data_col85[62] <= data_col85[61];
   data_col85[63] <= data_col85[62];
   data_col85[64] <= data_col85[63];
   data_col85[65] <= data_col85[64];
   data_col85[66] <= data_col85[65];
   data_col85[67] <= data_col85[66];
   data_col85[68] <= data_col85[67];
   data_col85[69] <= data_col85[68];
   data_col85[70] <= data_col85[69];
   data_col85[71] <= data_col85[70];
   data_col85[72] <= data_col85[71];
   data_col85[73] <= data_col85[72];
   data_col85[74] <= data_col85[73];
   data_col85[75] <= data_col85[74];
   data_col85[76] <= data_col85[75];
   data_col85[77] <= data_col85[76];
   data_col85[78] <= data_col85[77];
   data_col85[79] <= data_col85[78];
   data_col85[80] <= data_col85[79];
   data_col85[81] <= data_col85[80];
   data_col85[82] <= data_col85[81];
   data_col85[83] <= data_col85[82];
   data_col85[84] <= data_col85[83];
   data_col85[85] <= data_col85[84];

   data_col86[1] <= data[14];
   data_col86[2] <= data_col86[1];
   data_col86[3] <= data_col86[2];
   data_col86[4] <= data_col86[3];
   data_col86[5] <= data_col86[4];
   data_col86[6] <= data_col86[5];
   data_col86[7] <= data_col86[6];
   data_col86[8] <= data_col86[7];
   data_col86[9] <= data_col86[8];
   data_col86[10] <= data_col86[9];
   data_col86[11] <= data_col86[10];
   data_col86[12] <= data_col86[11];
   data_col86[13] <= data_col86[12];
   data_col86[14] <= data_col86[13];
   data_col86[15] <= data_col86[14];
   data_col86[16] <= data_col86[15];
   data_col86[17] <= data_col86[16];
   data_col86[18] <= data_col86[17];
   data_col86[19] <= data_col86[18];
   data_col86[20] <= data_col86[19];
   data_col86[21] <= data_col86[20];
   data_col86[22] <= data_col86[21];
   data_col86[23] <= data_col86[22];
   data_col86[24] <= data_col86[23];
   data_col86[25] <= data_col86[24];
   data_col86[26] <= data_col86[25];
   data_col86[27] <= data_col86[26];
   data_col86[28] <= data_col86[27];
   data_col86[29] <= data_col86[28];
   data_col86[30] <= data_col86[29];
   data_col86[31] <= data_col86[30];
   data_col86[32] <= data_col86[31];
   data_col86[33] <= data_col86[32];
   data_col86[34] <= data_col86[33];
   data_col86[35] <= data_col86[34];
   data_col86[36] <= data_col86[35];
   data_col86[37] <= data_col86[36];
   data_col86[38] <= data_col86[37];
   data_col86[39] <= data_col86[38];
   data_col86[40] <= data_col86[39];
   data_col86[41] <= data_col86[40];
   data_col86[42] <= data_col86[41];
   data_col86[43] <= data_col86[42];
   data_col86[44] <= data_col86[43];
   data_col86[45] <= data_col86[44];
   data_col86[46] <= data_col86[45];
   data_col86[47] <= data_col86[46];
   data_col86[48] <= data_col86[47];
   data_col86[49] <= data_col86[48];
   data_col86[50] <= data_col86[49];
   data_col86[51] <= data_col86[50];
   data_col86[52] <= data_col86[51];
   data_col86[53] <= data_col86[52];
   data_col86[54] <= data_col86[53];
   data_col86[55] <= data_col86[54];
   data_col86[56] <= data_col86[55];
   data_col86[57] <= data_col86[56];
   data_col86[58] <= data_col86[57];
   data_col86[59] <= data_col86[58];
   data_col86[60] <= data_col86[59];
   data_col86[61] <= data_col86[60];
   data_col86[62] <= data_col86[61];
   data_col86[63] <= data_col86[62];
   data_col86[64] <= data_col86[63];
   data_col86[65] <= data_col86[64];
   data_col86[66] <= data_col86[65];
   data_col86[67] <= data_col86[66];
   data_col86[68] <= data_col86[67];
   data_col86[69] <= data_col86[68];
   data_col86[70] <= data_col86[69];
   data_col86[71] <= data_col86[70];
   data_col86[72] <= data_col86[71];
   data_col86[73] <= data_col86[72];
   data_col86[74] <= data_col86[73];
   data_col86[75] <= data_col86[74];
   data_col86[76] <= data_col86[75];
   data_col86[77] <= data_col86[76];
   data_col86[78] <= data_col86[77];
   data_col86[79] <= data_col86[78];
   data_col86[80] <= data_col86[79];
   data_col86[81] <= data_col86[80];
   data_col86[82] <= data_col86[81];
   data_col86[83] <= data_col86[82];
   data_col86[84] <= data_col86[83];
   data_col86[85] <= data_col86[84];
   data_col86[86] <= data_col86[85];

   data_col87[1] <= data[13];
   data_col87[2] <= data_col87[1];
   data_col87[3] <= data_col87[2];
   data_col87[4] <= data_col87[3];
   data_col87[5] <= data_col87[4];
   data_col87[6] <= data_col87[5];
   data_col87[7] <= data_col87[6];
   data_col87[8] <= data_col87[7];
   data_col87[9] <= data_col87[8];
   data_col87[10] <= data_col87[9];
   data_col87[11] <= data_col87[10];
   data_col87[12] <= data_col87[11];
   data_col87[13] <= data_col87[12];
   data_col87[14] <= data_col87[13];
   data_col87[15] <= data_col87[14];
   data_col87[16] <= data_col87[15];
   data_col87[17] <= data_col87[16];
   data_col87[18] <= data_col87[17];
   data_col87[19] <= data_col87[18];
   data_col87[20] <= data_col87[19];
   data_col87[21] <= data_col87[20];
   data_col87[22] <= data_col87[21];
   data_col87[23] <= data_col87[22];
   data_col87[24] <= data_col87[23];
   data_col87[25] <= data_col87[24];
   data_col87[26] <= data_col87[25];
   data_col87[27] <= data_col87[26];
   data_col87[28] <= data_col87[27];
   data_col87[29] <= data_col87[28];
   data_col87[30] <= data_col87[29];
   data_col87[31] <= data_col87[30];
   data_col87[32] <= data_col87[31];
   data_col87[33] <= data_col87[32];
   data_col87[34] <= data_col87[33];
   data_col87[35] <= data_col87[34];
   data_col87[36] <= data_col87[35];
   data_col87[37] <= data_col87[36];
   data_col87[38] <= data_col87[37];
   data_col87[39] <= data_col87[38];
   data_col87[40] <= data_col87[39];
   data_col87[41] <= data_col87[40];
   data_col87[42] <= data_col87[41];
   data_col87[43] <= data_col87[42];
   data_col87[44] <= data_col87[43];
   data_col87[45] <= data_col87[44];
   data_col87[46] <= data_col87[45];
   data_col87[47] <= data_col87[46];
   data_col87[48] <= data_col87[47];
   data_col87[49] <= data_col87[48];
   data_col87[50] <= data_col87[49];
   data_col87[51] <= data_col87[50];
   data_col87[52] <= data_col87[51];
   data_col87[53] <= data_col87[52];
   data_col87[54] <= data_col87[53];
   data_col87[55] <= data_col87[54];
   data_col87[56] <= data_col87[55];
   data_col87[57] <= data_col87[56];
   data_col87[58] <= data_col87[57];
   data_col87[59] <= data_col87[58];
   data_col87[60] <= data_col87[59];
   data_col87[61] <= data_col87[60];
   data_col87[62] <= data_col87[61];
   data_col87[63] <= data_col87[62];
   data_col87[64] <= data_col87[63];
   data_col87[65] <= data_col87[64];
   data_col87[66] <= data_col87[65];
   data_col87[67] <= data_col87[66];
   data_col87[68] <= data_col87[67];
   data_col87[69] <= data_col87[68];
   data_col87[70] <= data_col87[69];
   data_col87[71] <= data_col87[70];
   data_col87[72] <= data_col87[71];
   data_col87[73] <= data_col87[72];
   data_col87[74] <= data_col87[73];
   data_col87[75] <= data_col87[74];
   data_col87[76] <= data_col87[75];
   data_col87[77] <= data_col87[76];
   data_col87[78] <= data_col87[77];
   data_col87[79] <= data_col87[78];
   data_col87[80] <= data_col87[79];
   data_col87[81] <= data_col87[80];
   data_col87[82] <= data_col87[81];
   data_col87[83] <= data_col87[82];
   data_col87[84] <= data_col87[83];
   data_col87[85] <= data_col87[84];
   data_col87[86] <= data_col87[85];
   data_col87[87] <= data_col87[86];

   data_col88[1] <= data[12];
   data_col88[2] <= data_col88[1];
   data_col88[3] <= data_col88[2];
   data_col88[4] <= data_col88[3];
   data_col88[5] <= data_col88[4];
   data_col88[6] <= data_col88[5];
   data_col88[7] <= data_col88[6];
   data_col88[8] <= data_col88[7];
   data_col88[9] <= data_col88[8];
   data_col88[10] <= data_col88[9];
   data_col88[11] <= data_col88[10];
   data_col88[12] <= data_col88[11];
   data_col88[13] <= data_col88[12];
   data_col88[14] <= data_col88[13];
   data_col88[15] <= data_col88[14];
   data_col88[16] <= data_col88[15];
   data_col88[17] <= data_col88[16];
   data_col88[18] <= data_col88[17];
   data_col88[19] <= data_col88[18];
   data_col88[20] <= data_col88[19];
   data_col88[21] <= data_col88[20];
   data_col88[22] <= data_col88[21];
   data_col88[23] <= data_col88[22];
   data_col88[24] <= data_col88[23];
   data_col88[25] <= data_col88[24];
   data_col88[26] <= data_col88[25];
   data_col88[27] <= data_col88[26];
   data_col88[28] <= data_col88[27];
   data_col88[29] <= data_col88[28];
   data_col88[30] <= data_col88[29];
   data_col88[31] <= data_col88[30];
   data_col88[32] <= data_col88[31];
   data_col88[33] <= data_col88[32];
   data_col88[34] <= data_col88[33];
   data_col88[35] <= data_col88[34];
   data_col88[36] <= data_col88[35];
   data_col88[37] <= data_col88[36];
   data_col88[38] <= data_col88[37];
   data_col88[39] <= data_col88[38];
   data_col88[40] <= data_col88[39];
   data_col88[41] <= data_col88[40];
   data_col88[42] <= data_col88[41];
   data_col88[43] <= data_col88[42];
   data_col88[44] <= data_col88[43];
   data_col88[45] <= data_col88[44];
   data_col88[46] <= data_col88[45];
   data_col88[47] <= data_col88[46];
   data_col88[48] <= data_col88[47];
   data_col88[49] <= data_col88[48];
   data_col88[50] <= data_col88[49];
   data_col88[51] <= data_col88[50];
   data_col88[52] <= data_col88[51];
   data_col88[53] <= data_col88[52];
   data_col88[54] <= data_col88[53];
   data_col88[55] <= data_col88[54];
   data_col88[56] <= data_col88[55];
   data_col88[57] <= data_col88[56];
   data_col88[58] <= data_col88[57];
   data_col88[59] <= data_col88[58];
   data_col88[60] <= data_col88[59];
   data_col88[61] <= data_col88[60];
   data_col88[62] <= data_col88[61];
   data_col88[63] <= data_col88[62];
   data_col88[64] <= data_col88[63];
   data_col88[65] <= data_col88[64];
   data_col88[66] <= data_col88[65];
   data_col88[67] <= data_col88[66];
   data_col88[68] <= data_col88[67];
   data_col88[69] <= data_col88[68];
   data_col88[70] <= data_col88[69];
   data_col88[71] <= data_col88[70];
   data_col88[72] <= data_col88[71];
   data_col88[73] <= data_col88[72];
   data_col88[74] <= data_col88[73];
   data_col88[75] <= data_col88[74];
   data_col88[76] <= data_col88[75];
   data_col88[77] <= data_col88[76];
   data_col88[78] <= data_col88[77];
   data_col88[79] <= data_col88[78];
   data_col88[80] <= data_col88[79];
   data_col88[81] <= data_col88[80];
   data_col88[82] <= data_col88[81];
   data_col88[83] <= data_col88[82];
   data_col88[84] <= data_col88[83];
   data_col88[85] <= data_col88[84];
   data_col88[86] <= data_col88[85];
   data_col88[87] <= data_col88[86];
   data_col88[88] <= data_col88[87];

   data_col89[1] <= data[11];
   data_col89[2] <= data_col89[1];
   data_col89[3] <= data_col89[2];
   data_col89[4] <= data_col89[3];
   data_col89[5] <= data_col89[4];
   data_col89[6] <= data_col89[5];
   data_col89[7] <= data_col89[6];
   data_col89[8] <= data_col89[7];
   data_col89[9] <= data_col89[8];
   data_col89[10] <= data_col89[9];
   data_col89[11] <= data_col89[10];
   data_col89[12] <= data_col89[11];
   data_col89[13] <= data_col89[12];
   data_col89[14] <= data_col89[13];
   data_col89[15] <= data_col89[14];
   data_col89[16] <= data_col89[15];
   data_col89[17] <= data_col89[16];
   data_col89[18] <= data_col89[17];
   data_col89[19] <= data_col89[18];
   data_col89[20] <= data_col89[19];
   data_col89[21] <= data_col89[20];
   data_col89[22] <= data_col89[21];
   data_col89[23] <= data_col89[22];
   data_col89[24] <= data_col89[23];
   data_col89[25] <= data_col89[24];
   data_col89[26] <= data_col89[25];
   data_col89[27] <= data_col89[26];
   data_col89[28] <= data_col89[27];
   data_col89[29] <= data_col89[28];
   data_col89[30] <= data_col89[29];
   data_col89[31] <= data_col89[30];
   data_col89[32] <= data_col89[31];
   data_col89[33] <= data_col89[32];
   data_col89[34] <= data_col89[33];
   data_col89[35] <= data_col89[34];
   data_col89[36] <= data_col89[35];
   data_col89[37] <= data_col89[36];
   data_col89[38] <= data_col89[37];
   data_col89[39] <= data_col89[38];
   data_col89[40] <= data_col89[39];
   data_col89[41] <= data_col89[40];
   data_col89[42] <= data_col89[41];
   data_col89[43] <= data_col89[42];
   data_col89[44] <= data_col89[43];
   data_col89[45] <= data_col89[44];
   data_col89[46] <= data_col89[45];
   data_col89[47] <= data_col89[46];
   data_col89[48] <= data_col89[47];
   data_col89[49] <= data_col89[48];
   data_col89[50] <= data_col89[49];
   data_col89[51] <= data_col89[50];
   data_col89[52] <= data_col89[51];
   data_col89[53] <= data_col89[52];
   data_col89[54] <= data_col89[53];
   data_col89[55] <= data_col89[54];
   data_col89[56] <= data_col89[55];
   data_col89[57] <= data_col89[56];
   data_col89[58] <= data_col89[57];
   data_col89[59] <= data_col89[58];
   data_col89[60] <= data_col89[59];
   data_col89[61] <= data_col89[60];
   data_col89[62] <= data_col89[61];
   data_col89[63] <= data_col89[62];
   data_col89[64] <= data_col89[63];
   data_col89[65] <= data_col89[64];
   data_col89[66] <= data_col89[65];
   data_col89[67] <= data_col89[66];
   data_col89[68] <= data_col89[67];
   data_col89[69] <= data_col89[68];
   data_col89[70] <= data_col89[69];
   data_col89[71] <= data_col89[70];
   data_col89[72] <= data_col89[71];
   data_col89[73] <= data_col89[72];
   data_col89[74] <= data_col89[73];
   data_col89[75] <= data_col89[74];
   data_col89[76] <= data_col89[75];
   data_col89[77] <= data_col89[76];
   data_col89[78] <= data_col89[77];
   data_col89[79] <= data_col89[78];
   data_col89[80] <= data_col89[79];
   data_col89[81] <= data_col89[80];
   data_col89[82] <= data_col89[81];
   data_col89[83] <= data_col89[82];
   data_col89[84] <= data_col89[83];
   data_col89[85] <= data_col89[84];
   data_col89[86] <= data_col89[85];
   data_col89[87] <= data_col89[86];
   data_col89[88] <= data_col89[87];
   data_col89[89] <= data_col89[88];

   data_col90[1] <= data[10];
   data_col90[2] <= data_col90[1];
   data_col90[3] <= data_col90[2];
   data_col90[4] <= data_col90[3];
   data_col90[5] <= data_col90[4];
   data_col90[6] <= data_col90[5];
   data_col90[7] <= data_col90[6];
   data_col90[8] <= data_col90[7];
   data_col90[9] <= data_col90[8];
   data_col90[10] <= data_col90[9];
   data_col90[11] <= data_col90[10];
   data_col90[12] <= data_col90[11];
   data_col90[13] <= data_col90[12];
   data_col90[14] <= data_col90[13];
   data_col90[15] <= data_col90[14];
   data_col90[16] <= data_col90[15];
   data_col90[17] <= data_col90[16];
   data_col90[18] <= data_col90[17];
   data_col90[19] <= data_col90[18];
   data_col90[20] <= data_col90[19];
   data_col90[21] <= data_col90[20];
   data_col90[22] <= data_col90[21];
   data_col90[23] <= data_col90[22];
   data_col90[24] <= data_col90[23];
   data_col90[25] <= data_col90[24];
   data_col90[26] <= data_col90[25];
   data_col90[27] <= data_col90[26];
   data_col90[28] <= data_col90[27];
   data_col90[29] <= data_col90[28];
   data_col90[30] <= data_col90[29];
   data_col90[31] <= data_col90[30];
   data_col90[32] <= data_col90[31];
   data_col90[33] <= data_col90[32];
   data_col90[34] <= data_col90[33];
   data_col90[35] <= data_col90[34];
   data_col90[36] <= data_col90[35];
   data_col90[37] <= data_col90[36];
   data_col90[38] <= data_col90[37];
   data_col90[39] <= data_col90[38];
   data_col90[40] <= data_col90[39];
   data_col90[41] <= data_col90[40];
   data_col90[42] <= data_col90[41];
   data_col90[43] <= data_col90[42];
   data_col90[44] <= data_col90[43];
   data_col90[45] <= data_col90[44];
   data_col90[46] <= data_col90[45];
   data_col90[47] <= data_col90[46];
   data_col90[48] <= data_col90[47];
   data_col90[49] <= data_col90[48];
   data_col90[50] <= data_col90[49];
   data_col90[51] <= data_col90[50];
   data_col90[52] <= data_col90[51];
   data_col90[53] <= data_col90[52];
   data_col90[54] <= data_col90[53];
   data_col90[55] <= data_col90[54];
   data_col90[56] <= data_col90[55];
   data_col90[57] <= data_col90[56];
   data_col90[58] <= data_col90[57];
   data_col90[59] <= data_col90[58];
   data_col90[60] <= data_col90[59];
   data_col90[61] <= data_col90[60];
   data_col90[62] <= data_col90[61];
   data_col90[63] <= data_col90[62];
   data_col90[64] <= data_col90[63];
   data_col90[65] <= data_col90[64];
   data_col90[66] <= data_col90[65];
   data_col90[67] <= data_col90[66];
   data_col90[68] <= data_col90[67];
   data_col90[69] <= data_col90[68];
   data_col90[70] <= data_col90[69];
   data_col90[71] <= data_col90[70];
   data_col90[72] <= data_col90[71];
   data_col90[73] <= data_col90[72];
   data_col90[74] <= data_col90[73];
   data_col90[75] <= data_col90[74];
   data_col90[76] <= data_col90[75];
   data_col90[77] <= data_col90[76];
   data_col90[78] <= data_col90[77];
   data_col90[79] <= data_col90[78];
   data_col90[80] <= data_col90[79];
   data_col90[81] <= data_col90[80];
   data_col90[82] <= data_col90[81];
   data_col90[83] <= data_col90[82];
   data_col90[84] <= data_col90[83];
   data_col90[85] <= data_col90[84];
   data_col90[86] <= data_col90[85];
   data_col90[87] <= data_col90[86];
   data_col90[88] <= data_col90[87];
   data_col90[89] <= data_col90[88];
   data_col90[90] <= data_col90[89];

   data_col91[1] <= data[9];
   data_col91[2] <= data_col91[1];
   data_col91[3] <= data_col91[2];
   data_col91[4] <= data_col91[3];
   data_col91[5] <= data_col91[4];
   data_col91[6] <= data_col91[5];
   data_col91[7] <= data_col91[6];
   data_col91[8] <= data_col91[7];
   data_col91[9] <= data_col91[8];
   data_col91[10] <= data_col91[9];
   data_col91[11] <= data_col91[10];
   data_col91[12] <= data_col91[11];
   data_col91[13] <= data_col91[12];
   data_col91[14] <= data_col91[13];
   data_col91[15] <= data_col91[14];
   data_col91[16] <= data_col91[15];
   data_col91[17] <= data_col91[16];
   data_col91[18] <= data_col91[17];
   data_col91[19] <= data_col91[18];
   data_col91[20] <= data_col91[19];
   data_col91[21] <= data_col91[20];
   data_col91[22] <= data_col91[21];
   data_col91[23] <= data_col91[22];
   data_col91[24] <= data_col91[23];
   data_col91[25] <= data_col91[24];
   data_col91[26] <= data_col91[25];
   data_col91[27] <= data_col91[26];
   data_col91[28] <= data_col91[27];
   data_col91[29] <= data_col91[28];
   data_col91[30] <= data_col91[29];
   data_col91[31] <= data_col91[30];
   data_col91[32] <= data_col91[31];
   data_col91[33] <= data_col91[32];
   data_col91[34] <= data_col91[33];
   data_col91[35] <= data_col91[34];
   data_col91[36] <= data_col91[35];
   data_col91[37] <= data_col91[36];
   data_col91[38] <= data_col91[37];
   data_col91[39] <= data_col91[38];
   data_col91[40] <= data_col91[39];
   data_col91[41] <= data_col91[40];
   data_col91[42] <= data_col91[41];
   data_col91[43] <= data_col91[42];
   data_col91[44] <= data_col91[43];
   data_col91[45] <= data_col91[44];
   data_col91[46] <= data_col91[45];
   data_col91[47] <= data_col91[46];
   data_col91[48] <= data_col91[47];
   data_col91[49] <= data_col91[48];
   data_col91[50] <= data_col91[49];
   data_col91[51] <= data_col91[50];
   data_col91[52] <= data_col91[51];
   data_col91[53] <= data_col91[52];
   data_col91[54] <= data_col91[53];
   data_col91[55] <= data_col91[54];
   data_col91[56] <= data_col91[55];
   data_col91[57] <= data_col91[56];
   data_col91[58] <= data_col91[57];
   data_col91[59] <= data_col91[58];
   data_col91[60] <= data_col91[59];
   data_col91[61] <= data_col91[60];
   data_col91[62] <= data_col91[61];
   data_col91[63] <= data_col91[62];
   data_col91[64] <= data_col91[63];
   data_col91[65] <= data_col91[64];
   data_col91[66] <= data_col91[65];
   data_col91[67] <= data_col91[66];
   data_col91[68] <= data_col91[67];
   data_col91[69] <= data_col91[68];
   data_col91[70] <= data_col91[69];
   data_col91[71] <= data_col91[70];
   data_col91[72] <= data_col91[71];
   data_col91[73] <= data_col91[72];
   data_col91[74] <= data_col91[73];
   data_col91[75] <= data_col91[74];
   data_col91[76] <= data_col91[75];
   data_col91[77] <= data_col91[76];
   data_col91[78] <= data_col91[77];
   data_col91[79] <= data_col91[78];
   data_col91[80] <= data_col91[79];
   data_col91[81] <= data_col91[80];
   data_col91[82] <= data_col91[81];
   data_col91[83] <= data_col91[82];
   data_col91[84] <= data_col91[83];
   data_col91[85] <= data_col91[84];
   data_col91[86] <= data_col91[85];
   data_col91[87] <= data_col91[86];
   data_col91[88] <= data_col91[87];
   data_col91[89] <= data_col91[88];
   data_col91[90] <= data_col91[89];
   data_col91[91] <= data_col91[90];

   data_col92[1] <= data[8];
   data_col92[2] <= data_col92[1];
   data_col92[3] <= data_col92[2];
   data_col92[4] <= data_col92[3];
   data_col92[5] <= data_col92[4];
   data_col92[6] <= data_col92[5];
   data_col92[7] <= data_col92[6];
   data_col92[8] <= data_col92[7];
   data_col92[9] <= data_col92[8];
   data_col92[10] <= data_col92[9];
   data_col92[11] <= data_col92[10];
   data_col92[12] <= data_col92[11];
   data_col92[13] <= data_col92[12];
   data_col92[14] <= data_col92[13];
   data_col92[15] <= data_col92[14];
   data_col92[16] <= data_col92[15];
   data_col92[17] <= data_col92[16];
   data_col92[18] <= data_col92[17];
   data_col92[19] <= data_col92[18];
   data_col92[20] <= data_col92[19];
   data_col92[21] <= data_col92[20];
   data_col92[22] <= data_col92[21];
   data_col92[23] <= data_col92[22];
   data_col92[24] <= data_col92[23];
   data_col92[25] <= data_col92[24];
   data_col92[26] <= data_col92[25];
   data_col92[27] <= data_col92[26];
   data_col92[28] <= data_col92[27];
   data_col92[29] <= data_col92[28];
   data_col92[30] <= data_col92[29];
   data_col92[31] <= data_col92[30];
   data_col92[32] <= data_col92[31];
   data_col92[33] <= data_col92[32];
   data_col92[34] <= data_col92[33];
   data_col92[35] <= data_col92[34];
   data_col92[36] <= data_col92[35];
   data_col92[37] <= data_col92[36];
   data_col92[38] <= data_col92[37];
   data_col92[39] <= data_col92[38];
   data_col92[40] <= data_col92[39];
   data_col92[41] <= data_col92[40];
   data_col92[42] <= data_col92[41];
   data_col92[43] <= data_col92[42];
   data_col92[44] <= data_col92[43];
   data_col92[45] <= data_col92[44];
   data_col92[46] <= data_col92[45];
   data_col92[47] <= data_col92[46];
   data_col92[48] <= data_col92[47];
   data_col92[49] <= data_col92[48];
   data_col92[50] <= data_col92[49];
   data_col92[51] <= data_col92[50];
   data_col92[52] <= data_col92[51];
   data_col92[53] <= data_col92[52];
   data_col92[54] <= data_col92[53];
   data_col92[55] <= data_col92[54];
   data_col92[56] <= data_col92[55];
   data_col92[57] <= data_col92[56];
   data_col92[58] <= data_col92[57];
   data_col92[59] <= data_col92[58];
   data_col92[60] <= data_col92[59];
   data_col92[61] <= data_col92[60];
   data_col92[62] <= data_col92[61];
   data_col92[63] <= data_col92[62];
   data_col92[64] <= data_col92[63];
   data_col92[65] <= data_col92[64];
   data_col92[66] <= data_col92[65];
   data_col92[67] <= data_col92[66];
   data_col92[68] <= data_col92[67];
   data_col92[69] <= data_col92[68];
   data_col92[70] <= data_col92[69];
   data_col92[71] <= data_col92[70];
   data_col92[72] <= data_col92[71];
   data_col92[73] <= data_col92[72];
   data_col92[74] <= data_col92[73];
   data_col92[75] <= data_col92[74];
   data_col92[76] <= data_col92[75];
   data_col92[77] <= data_col92[76];
   data_col92[78] <= data_col92[77];
   data_col92[79] <= data_col92[78];
   data_col92[80] <= data_col92[79];
   data_col92[81] <= data_col92[80];
   data_col92[82] <= data_col92[81];
   data_col92[83] <= data_col92[82];
   data_col92[84] <= data_col92[83];
   data_col92[85] <= data_col92[84];
   data_col92[86] <= data_col92[85];
   data_col92[87] <= data_col92[86];
   data_col92[88] <= data_col92[87];
   data_col92[89] <= data_col92[88];
   data_col92[90] <= data_col92[89];
   data_col92[91] <= data_col92[90];
   data_col92[92] <= data_col92[91];

   data_col93[1] <= data[7];
   data_col93[2] <= data_col93[1];
   data_col93[3] <= data_col93[2];
   data_col93[4] <= data_col93[3];
   data_col93[5] <= data_col93[4];
   data_col93[6] <= data_col93[5];
   data_col93[7] <= data_col93[6];
   data_col93[8] <= data_col93[7];
   data_col93[9] <= data_col93[8];
   data_col93[10] <= data_col93[9];
   data_col93[11] <= data_col93[10];
   data_col93[12] <= data_col93[11];
   data_col93[13] <= data_col93[12];
   data_col93[14] <= data_col93[13];
   data_col93[15] <= data_col93[14];
   data_col93[16] <= data_col93[15];
   data_col93[17] <= data_col93[16];
   data_col93[18] <= data_col93[17];
   data_col93[19] <= data_col93[18];
   data_col93[20] <= data_col93[19];
   data_col93[21] <= data_col93[20];
   data_col93[22] <= data_col93[21];
   data_col93[23] <= data_col93[22];
   data_col93[24] <= data_col93[23];
   data_col93[25] <= data_col93[24];
   data_col93[26] <= data_col93[25];
   data_col93[27] <= data_col93[26];
   data_col93[28] <= data_col93[27];
   data_col93[29] <= data_col93[28];
   data_col93[30] <= data_col93[29];
   data_col93[31] <= data_col93[30];
   data_col93[32] <= data_col93[31];
   data_col93[33] <= data_col93[32];
   data_col93[34] <= data_col93[33];
   data_col93[35] <= data_col93[34];
   data_col93[36] <= data_col93[35];
   data_col93[37] <= data_col93[36];
   data_col93[38] <= data_col93[37];
   data_col93[39] <= data_col93[38];
   data_col93[40] <= data_col93[39];
   data_col93[41] <= data_col93[40];
   data_col93[42] <= data_col93[41];
   data_col93[43] <= data_col93[42];
   data_col93[44] <= data_col93[43];
   data_col93[45] <= data_col93[44];
   data_col93[46] <= data_col93[45];
   data_col93[47] <= data_col93[46];
   data_col93[48] <= data_col93[47];
   data_col93[49] <= data_col93[48];
   data_col93[50] <= data_col93[49];
   data_col93[51] <= data_col93[50];
   data_col93[52] <= data_col93[51];
   data_col93[53] <= data_col93[52];
   data_col93[54] <= data_col93[53];
   data_col93[55] <= data_col93[54];
   data_col93[56] <= data_col93[55];
   data_col93[57] <= data_col93[56];
   data_col93[58] <= data_col93[57];
   data_col93[59] <= data_col93[58];
   data_col93[60] <= data_col93[59];
   data_col93[61] <= data_col93[60];
   data_col93[62] <= data_col93[61];
   data_col93[63] <= data_col93[62];
   data_col93[64] <= data_col93[63];
   data_col93[65] <= data_col93[64];
   data_col93[66] <= data_col93[65];
   data_col93[67] <= data_col93[66];
   data_col93[68] <= data_col93[67];
   data_col93[69] <= data_col93[68];
   data_col93[70] <= data_col93[69];
   data_col93[71] <= data_col93[70];
   data_col93[72] <= data_col93[71];
   data_col93[73] <= data_col93[72];
   data_col93[74] <= data_col93[73];
   data_col93[75] <= data_col93[74];
   data_col93[76] <= data_col93[75];
   data_col93[77] <= data_col93[76];
   data_col93[78] <= data_col93[77];
   data_col93[79] <= data_col93[78];
   data_col93[80] <= data_col93[79];
   data_col93[81] <= data_col93[80];
   data_col93[82] <= data_col93[81];
   data_col93[83] <= data_col93[82];
   data_col93[84] <= data_col93[83];
   data_col93[85] <= data_col93[84];
   data_col93[86] <= data_col93[85];
   data_col93[87] <= data_col93[86];
   data_col93[88] <= data_col93[87];
   data_col93[89] <= data_col93[88];
   data_col93[90] <= data_col93[89];
   data_col93[91] <= data_col93[90];
   data_col93[92] <= data_col93[91];
   data_col93[93] <= data_col93[92];

   data_col94[1] <= data[6];
   data_col94[2] <= data_col94[1];
   data_col94[3] <= data_col94[2];
   data_col94[4] <= data_col94[3];
   data_col94[5] <= data_col94[4];
   data_col94[6] <= data_col94[5];
   data_col94[7] <= data_col94[6];
   data_col94[8] <= data_col94[7];
   data_col94[9] <= data_col94[8];
   data_col94[10] <= data_col94[9];
   data_col94[11] <= data_col94[10];
   data_col94[12] <= data_col94[11];
   data_col94[13] <= data_col94[12];
   data_col94[14] <= data_col94[13];
   data_col94[15] <= data_col94[14];
   data_col94[16] <= data_col94[15];
   data_col94[17] <= data_col94[16];
   data_col94[18] <= data_col94[17];
   data_col94[19] <= data_col94[18];
   data_col94[20] <= data_col94[19];
   data_col94[21] <= data_col94[20];
   data_col94[22] <= data_col94[21];
   data_col94[23] <= data_col94[22];
   data_col94[24] <= data_col94[23];
   data_col94[25] <= data_col94[24];
   data_col94[26] <= data_col94[25];
   data_col94[27] <= data_col94[26];
   data_col94[28] <= data_col94[27];
   data_col94[29] <= data_col94[28];
   data_col94[30] <= data_col94[29];
   data_col94[31] <= data_col94[30];
   data_col94[32] <= data_col94[31];
   data_col94[33] <= data_col94[32];
   data_col94[34] <= data_col94[33];
   data_col94[35] <= data_col94[34];
   data_col94[36] <= data_col94[35];
   data_col94[37] <= data_col94[36];
   data_col94[38] <= data_col94[37];
   data_col94[39] <= data_col94[38];
   data_col94[40] <= data_col94[39];
   data_col94[41] <= data_col94[40];
   data_col94[42] <= data_col94[41];
   data_col94[43] <= data_col94[42];
   data_col94[44] <= data_col94[43];
   data_col94[45] <= data_col94[44];
   data_col94[46] <= data_col94[45];
   data_col94[47] <= data_col94[46];
   data_col94[48] <= data_col94[47];
   data_col94[49] <= data_col94[48];
   data_col94[50] <= data_col94[49];
   data_col94[51] <= data_col94[50];
   data_col94[52] <= data_col94[51];
   data_col94[53] <= data_col94[52];
   data_col94[54] <= data_col94[53];
   data_col94[55] <= data_col94[54];
   data_col94[56] <= data_col94[55];
   data_col94[57] <= data_col94[56];
   data_col94[58] <= data_col94[57];
   data_col94[59] <= data_col94[58];
   data_col94[60] <= data_col94[59];
   data_col94[61] <= data_col94[60];
   data_col94[62] <= data_col94[61];
   data_col94[63] <= data_col94[62];
   data_col94[64] <= data_col94[63];
   data_col94[65] <= data_col94[64];
   data_col94[66] <= data_col94[65];
   data_col94[67] <= data_col94[66];
   data_col94[68] <= data_col94[67];
   data_col94[69] <= data_col94[68];
   data_col94[70] <= data_col94[69];
   data_col94[71] <= data_col94[70];
   data_col94[72] <= data_col94[71];
   data_col94[73] <= data_col94[72];
   data_col94[74] <= data_col94[73];
   data_col94[75] <= data_col94[74];
   data_col94[76] <= data_col94[75];
   data_col94[77] <= data_col94[76];
   data_col94[78] <= data_col94[77];
   data_col94[79] <= data_col94[78];
   data_col94[80] <= data_col94[79];
   data_col94[81] <= data_col94[80];
   data_col94[82] <= data_col94[81];
   data_col94[83] <= data_col94[82];
   data_col94[84] <= data_col94[83];
   data_col94[85] <= data_col94[84];
   data_col94[86] <= data_col94[85];
   data_col94[87] <= data_col94[86];
   data_col94[88] <= data_col94[87];
   data_col94[89] <= data_col94[88];
   data_col94[90] <= data_col94[89];
   data_col94[91] <= data_col94[90];
   data_col94[92] <= data_col94[91];
   data_col94[93] <= data_col94[92];
   data_col94[94] <= data_col94[93];

   data_col95[1] <= data[5];
   data_col95[2] <= data_col95[1];
   data_col95[3] <= data_col95[2];
   data_col95[4] <= data_col95[3];
   data_col95[5] <= data_col95[4];
   data_col95[6] <= data_col95[5];
   data_col95[7] <= data_col95[6];
   data_col95[8] <= data_col95[7];
   data_col95[9] <= data_col95[8];
   data_col95[10] <= data_col95[9];
   data_col95[11] <= data_col95[10];
   data_col95[12] <= data_col95[11];
   data_col95[13] <= data_col95[12];
   data_col95[14] <= data_col95[13];
   data_col95[15] <= data_col95[14];
   data_col95[16] <= data_col95[15];
   data_col95[17] <= data_col95[16];
   data_col95[18] <= data_col95[17];
   data_col95[19] <= data_col95[18];
   data_col95[20] <= data_col95[19];
   data_col95[21] <= data_col95[20];
   data_col95[22] <= data_col95[21];
   data_col95[23] <= data_col95[22];
   data_col95[24] <= data_col95[23];
   data_col95[25] <= data_col95[24];
   data_col95[26] <= data_col95[25];
   data_col95[27] <= data_col95[26];
   data_col95[28] <= data_col95[27];
   data_col95[29] <= data_col95[28];
   data_col95[30] <= data_col95[29];
   data_col95[31] <= data_col95[30];
   data_col95[32] <= data_col95[31];
   data_col95[33] <= data_col95[32];
   data_col95[34] <= data_col95[33];
   data_col95[35] <= data_col95[34];
   data_col95[36] <= data_col95[35];
   data_col95[37] <= data_col95[36];
   data_col95[38] <= data_col95[37];
   data_col95[39] <= data_col95[38];
   data_col95[40] <= data_col95[39];
   data_col95[41] <= data_col95[40];
   data_col95[42] <= data_col95[41];
   data_col95[43] <= data_col95[42];
   data_col95[44] <= data_col95[43];
   data_col95[45] <= data_col95[44];
   data_col95[46] <= data_col95[45];
   data_col95[47] <= data_col95[46];
   data_col95[48] <= data_col95[47];
   data_col95[49] <= data_col95[48];
   data_col95[50] <= data_col95[49];
   data_col95[51] <= data_col95[50];
   data_col95[52] <= data_col95[51];
   data_col95[53] <= data_col95[52];
   data_col95[54] <= data_col95[53];
   data_col95[55] <= data_col95[54];
   data_col95[56] <= data_col95[55];
   data_col95[57] <= data_col95[56];
   data_col95[58] <= data_col95[57];
   data_col95[59] <= data_col95[58];
   data_col95[60] <= data_col95[59];
   data_col95[61] <= data_col95[60];
   data_col95[62] <= data_col95[61];
   data_col95[63] <= data_col95[62];
   data_col95[64] <= data_col95[63];
   data_col95[65] <= data_col95[64];
   data_col95[66] <= data_col95[65];
   data_col95[67] <= data_col95[66];
   data_col95[68] <= data_col95[67];
   data_col95[69] <= data_col95[68];
   data_col95[70] <= data_col95[69];
   data_col95[71] <= data_col95[70];
   data_col95[72] <= data_col95[71];
   data_col95[73] <= data_col95[72];
   data_col95[74] <= data_col95[73];
   data_col95[75] <= data_col95[74];
   data_col95[76] <= data_col95[75];
   data_col95[77] <= data_col95[76];
   data_col95[78] <= data_col95[77];
   data_col95[79] <= data_col95[78];
   data_col95[80] <= data_col95[79];
   data_col95[81] <= data_col95[80];
   data_col95[82] <= data_col95[81];
   data_col95[83] <= data_col95[82];
   data_col95[84] <= data_col95[83];
   data_col95[85] <= data_col95[84];
   data_col95[86] <= data_col95[85];
   data_col95[87] <= data_col95[86];
   data_col95[88] <= data_col95[87];
   data_col95[89] <= data_col95[88];
   data_col95[90] <= data_col95[89];
   data_col95[91] <= data_col95[90];
   data_col95[92] <= data_col95[91];
   data_col95[93] <= data_col95[92];
   data_col95[94] <= data_col95[93];
   data_col95[95] <= data_col95[94];

   data_col96[1] <= data[4];
   data_col96[2] <= data_col96[1];
   data_col96[3] <= data_col96[2];
   data_col96[4] <= data_col96[3];
   data_col96[5] <= data_col96[4];
   data_col96[6] <= data_col96[5];
   data_col96[7] <= data_col96[6];
   data_col96[8] <= data_col96[7];
   data_col96[9] <= data_col96[8];
   data_col96[10] <= data_col96[9];
   data_col96[11] <= data_col96[10];
   data_col96[12] <= data_col96[11];
   data_col96[13] <= data_col96[12];
   data_col96[14] <= data_col96[13];
   data_col96[15] <= data_col96[14];
   data_col96[16] <= data_col96[15];
   data_col96[17] <= data_col96[16];
   data_col96[18] <= data_col96[17];
   data_col96[19] <= data_col96[18];
   data_col96[20] <= data_col96[19];
   data_col96[21] <= data_col96[20];
   data_col96[22] <= data_col96[21];
   data_col96[23] <= data_col96[22];
   data_col96[24] <= data_col96[23];
   data_col96[25] <= data_col96[24];
   data_col96[26] <= data_col96[25];
   data_col96[27] <= data_col96[26];
   data_col96[28] <= data_col96[27];
   data_col96[29] <= data_col96[28];
   data_col96[30] <= data_col96[29];
   data_col96[31] <= data_col96[30];
   data_col96[32] <= data_col96[31];
   data_col96[33] <= data_col96[32];
   data_col96[34] <= data_col96[33];
   data_col96[35] <= data_col96[34];
   data_col96[36] <= data_col96[35];
   data_col96[37] <= data_col96[36];
   data_col96[38] <= data_col96[37];
   data_col96[39] <= data_col96[38];
   data_col96[40] <= data_col96[39];
   data_col96[41] <= data_col96[40];
   data_col96[42] <= data_col96[41];
   data_col96[43] <= data_col96[42];
   data_col96[44] <= data_col96[43];
   data_col96[45] <= data_col96[44];
   data_col96[46] <= data_col96[45];
   data_col96[47] <= data_col96[46];
   data_col96[48] <= data_col96[47];
   data_col96[49] <= data_col96[48];
   data_col96[50] <= data_col96[49];
   data_col96[51] <= data_col96[50];
   data_col96[52] <= data_col96[51];
   data_col96[53] <= data_col96[52];
   data_col96[54] <= data_col96[53];
   data_col96[55] <= data_col96[54];
   data_col96[56] <= data_col96[55];
   data_col96[57] <= data_col96[56];
   data_col96[58] <= data_col96[57];
   data_col96[59] <= data_col96[58];
   data_col96[60] <= data_col96[59];
   data_col96[61] <= data_col96[60];
   data_col96[62] <= data_col96[61];
   data_col96[63] <= data_col96[62];
   data_col96[64] <= data_col96[63];
   data_col96[65] <= data_col96[64];
   data_col96[66] <= data_col96[65];
   data_col96[67] <= data_col96[66];
   data_col96[68] <= data_col96[67];
   data_col96[69] <= data_col96[68];
   data_col96[70] <= data_col96[69];
   data_col96[71] <= data_col96[70];
   data_col96[72] <= data_col96[71];
   data_col96[73] <= data_col96[72];
   data_col96[74] <= data_col96[73];
   data_col96[75] <= data_col96[74];
   data_col96[76] <= data_col96[75];
   data_col96[77] <= data_col96[76];
   data_col96[78] <= data_col96[77];
   data_col96[79] <= data_col96[78];
   data_col96[80] <= data_col96[79];
   data_col96[81] <= data_col96[80];
   data_col96[82] <= data_col96[81];
   data_col96[83] <= data_col96[82];
   data_col96[84] <= data_col96[83];
   data_col96[85] <= data_col96[84];
   data_col96[86] <= data_col96[85];
   data_col96[87] <= data_col96[86];
   data_col96[88] <= data_col96[87];
   data_col96[89] <= data_col96[88];
   data_col96[90] <= data_col96[89];
   data_col96[91] <= data_col96[90];
   data_col96[92] <= data_col96[91];
   data_col96[93] <= data_col96[92];
   data_col96[94] <= data_col96[93];
   data_col96[95] <= data_col96[94];
   data_col96[96] <= data_col96[95];

   data_col97[1] <= data[3];
   data_col97[2] <= data_col97[1];
   data_col97[3] <= data_col97[2];
   data_col97[4] <= data_col97[3];
   data_col97[5] <= data_col97[4];
   data_col97[6] <= data_col97[5];
   data_col97[7] <= data_col97[6];
   data_col97[8] <= data_col97[7];
   data_col97[9] <= data_col97[8];
   data_col97[10] <= data_col97[9];
   data_col97[11] <= data_col97[10];
   data_col97[12] <= data_col97[11];
   data_col97[13] <= data_col97[12];
   data_col97[14] <= data_col97[13];
   data_col97[15] <= data_col97[14];
   data_col97[16] <= data_col97[15];
   data_col97[17] <= data_col97[16];
   data_col97[18] <= data_col97[17];
   data_col97[19] <= data_col97[18];
   data_col97[20] <= data_col97[19];
   data_col97[21] <= data_col97[20];
   data_col97[22] <= data_col97[21];
   data_col97[23] <= data_col97[22];
   data_col97[24] <= data_col97[23];
   data_col97[25] <= data_col97[24];
   data_col97[26] <= data_col97[25];
   data_col97[27] <= data_col97[26];
   data_col97[28] <= data_col97[27];
   data_col97[29] <= data_col97[28];
   data_col97[30] <= data_col97[29];
   data_col97[31] <= data_col97[30];
   data_col97[32] <= data_col97[31];
   data_col97[33] <= data_col97[32];
   data_col97[34] <= data_col97[33];
   data_col97[35] <= data_col97[34];
   data_col97[36] <= data_col97[35];
   data_col97[37] <= data_col97[36];
   data_col97[38] <= data_col97[37];
   data_col97[39] <= data_col97[38];
   data_col97[40] <= data_col97[39];
   data_col97[41] <= data_col97[40];
   data_col97[42] <= data_col97[41];
   data_col97[43] <= data_col97[42];
   data_col97[44] <= data_col97[43];
   data_col97[45] <= data_col97[44];
   data_col97[46] <= data_col97[45];
   data_col97[47] <= data_col97[46];
   data_col97[48] <= data_col97[47];
   data_col97[49] <= data_col97[48];
   data_col97[50] <= data_col97[49];
   data_col97[51] <= data_col97[50];
   data_col97[52] <= data_col97[51];
   data_col97[53] <= data_col97[52];
   data_col97[54] <= data_col97[53];
   data_col97[55] <= data_col97[54];
   data_col97[56] <= data_col97[55];
   data_col97[57] <= data_col97[56];
   data_col97[58] <= data_col97[57];
   data_col97[59] <= data_col97[58];
   data_col97[60] <= data_col97[59];
   data_col97[61] <= data_col97[60];
   data_col97[62] <= data_col97[61];
   data_col97[63] <= data_col97[62];
   data_col97[64] <= data_col97[63];
   data_col97[65] <= data_col97[64];
   data_col97[66] <= data_col97[65];
   data_col97[67] <= data_col97[66];
   data_col97[68] <= data_col97[67];
   data_col97[69] <= data_col97[68];
   data_col97[70] <= data_col97[69];
   data_col97[71] <= data_col97[70];
   data_col97[72] <= data_col97[71];
   data_col97[73] <= data_col97[72];
   data_col97[74] <= data_col97[73];
   data_col97[75] <= data_col97[74];
   data_col97[76] <= data_col97[75];
   data_col97[77] <= data_col97[76];
   data_col97[78] <= data_col97[77];
   data_col97[79] <= data_col97[78];
   data_col97[80] <= data_col97[79];
   data_col97[81] <= data_col97[80];
   data_col97[82] <= data_col97[81];
   data_col97[83] <= data_col97[82];
   data_col97[84] <= data_col97[83];
   data_col97[85] <= data_col97[84];
   data_col97[86] <= data_col97[85];
   data_col97[87] <= data_col97[86];
   data_col97[88] <= data_col97[87];
   data_col97[89] <= data_col97[88];
   data_col97[90] <= data_col97[89];
   data_col97[91] <= data_col97[90];
   data_col97[92] <= data_col97[91];
   data_col97[93] <= data_col97[92];
   data_col97[94] <= data_col97[93];
   data_col97[95] <= data_col97[94];
   data_col97[96] <= data_col97[95];
   data_col97[97] <= data_col97[96];

   data_col98[1] <= data[2];
   data_col98[2] <= data_col98[1];
   data_col98[3] <= data_col98[2];
   data_col98[4] <= data_col98[3];
   data_col98[5] <= data_col98[4];
   data_col98[6] <= data_col98[5];
   data_col98[7] <= data_col98[6];
   data_col98[8] <= data_col98[7];
   data_col98[9] <= data_col98[8];
   data_col98[10] <= data_col98[9];
   data_col98[11] <= data_col98[10];
   data_col98[12] <= data_col98[11];
   data_col98[13] <= data_col98[12];
   data_col98[14] <= data_col98[13];
   data_col98[15] <= data_col98[14];
   data_col98[16] <= data_col98[15];
   data_col98[17] <= data_col98[16];
   data_col98[18] <= data_col98[17];
   data_col98[19] <= data_col98[18];
   data_col98[20] <= data_col98[19];
   data_col98[21] <= data_col98[20];
   data_col98[22] <= data_col98[21];
   data_col98[23] <= data_col98[22];
   data_col98[24] <= data_col98[23];
   data_col98[25] <= data_col98[24];
   data_col98[26] <= data_col98[25];
   data_col98[27] <= data_col98[26];
   data_col98[28] <= data_col98[27];
   data_col98[29] <= data_col98[28];
   data_col98[30] <= data_col98[29];
   data_col98[31] <= data_col98[30];
   data_col98[32] <= data_col98[31];
   data_col98[33] <= data_col98[32];
   data_col98[34] <= data_col98[33];
   data_col98[35] <= data_col98[34];
   data_col98[36] <= data_col98[35];
   data_col98[37] <= data_col98[36];
   data_col98[38] <= data_col98[37];
   data_col98[39] <= data_col98[38];
   data_col98[40] <= data_col98[39];
   data_col98[41] <= data_col98[40];
   data_col98[42] <= data_col98[41];
   data_col98[43] <= data_col98[42];
   data_col98[44] <= data_col98[43];
   data_col98[45] <= data_col98[44];
   data_col98[46] <= data_col98[45];
   data_col98[47] <= data_col98[46];
   data_col98[48] <= data_col98[47];
   data_col98[49] <= data_col98[48];
   data_col98[50] <= data_col98[49];
   data_col98[51] <= data_col98[50];
   data_col98[52] <= data_col98[51];
   data_col98[53] <= data_col98[52];
   data_col98[54] <= data_col98[53];
   data_col98[55] <= data_col98[54];
   data_col98[56] <= data_col98[55];
   data_col98[57] <= data_col98[56];
   data_col98[58] <= data_col98[57];
   data_col98[59] <= data_col98[58];
   data_col98[60] <= data_col98[59];
   data_col98[61] <= data_col98[60];
   data_col98[62] <= data_col98[61];
   data_col98[63] <= data_col98[62];
   data_col98[64] <= data_col98[63];
   data_col98[65] <= data_col98[64];
   data_col98[66] <= data_col98[65];
   data_col98[67] <= data_col98[66];
   data_col98[68] <= data_col98[67];
   data_col98[69] <= data_col98[68];
   data_col98[70] <= data_col98[69];
   data_col98[71] <= data_col98[70];
   data_col98[72] <= data_col98[71];
   data_col98[73] <= data_col98[72];
   data_col98[74] <= data_col98[73];
   data_col98[75] <= data_col98[74];
   data_col98[76] <= data_col98[75];
   data_col98[77] <= data_col98[76];
   data_col98[78] <= data_col98[77];
   data_col98[79] <= data_col98[78];
   data_col98[80] <= data_col98[79];
   data_col98[81] <= data_col98[80];
   data_col98[82] <= data_col98[81];
   data_col98[83] <= data_col98[82];
   data_col98[84] <= data_col98[83];
   data_col98[85] <= data_col98[84];
   data_col98[86] <= data_col98[85];
   data_col98[87] <= data_col98[86];
   data_col98[88] <= data_col98[87];
   data_col98[89] <= data_col98[88];
   data_col98[90] <= data_col98[89];
   data_col98[91] <= data_col98[90];
   data_col98[92] <= data_col98[91];
   data_col98[93] <= data_col98[92];
   data_col98[94] <= data_col98[93];
   data_col98[95] <= data_col98[94];
   data_col98[96] <= data_col98[95];
   data_col98[97] <= data_col98[96];
   data_col98[98] <= data_col98[97];

   data_col99[1] <= data[1];
   data_col99[2] <= data_col99[1];
   data_col99[3] <= data_col99[2];
   data_col99[4] <= data_col99[3];
   data_col99[5] <= data_col99[4];
   data_col99[6] <= data_col99[5];
   data_col99[7] <= data_col99[6];
   data_col99[8] <= data_col99[7];
   data_col99[9] <= data_col99[8];
   data_col99[10] <= data_col99[9];
   data_col99[11] <= data_col99[10];
   data_col99[12] <= data_col99[11];
   data_col99[13] <= data_col99[12];
   data_col99[14] <= data_col99[13];
   data_col99[15] <= data_col99[14];
   data_col99[16] <= data_col99[15];
   data_col99[17] <= data_col99[16];
   data_col99[18] <= data_col99[17];
   data_col99[19] <= data_col99[18];
   data_col99[20] <= data_col99[19];
   data_col99[21] <= data_col99[20];
   data_col99[22] <= data_col99[21];
   data_col99[23] <= data_col99[22];
   data_col99[24] <= data_col99[23];
   data_col99[25] <= data_col99[24];
   data_col99[26] <= data_col99[25];
   data_col99[27] <= data_col99[26];
   data_col99[28] <= data_col99[27];
   data_col99[29] <= data_col99[28];
   data_col99[30] <= data_col99[29];
   data_col99[31] <= data_col99[30];
   data_col99[32] <= data_col99[31];
   data_col99[33] <= data_col99[32];
   data_col99[34] <= data_col99[33];
   data_col99[35] <= data_col99[34];
   data_col99[36] <= data_col99[35];
   data_col99[37] <= data_col99[36];
   data_col99[38] <= data_col99[37];
   data_col99[39] <= data_col99[38];
   data_col99[40] <= data_col99[39];
   data_col99[41] <= data_col99[40];
   data_col99[42] <= data_col99[41];
   data_col99[43] <= data_col99[42];
   data_col99[44] <= data_col99[43];
   data_col99[45] <= data_col99[44];
   data_col99[46] <= data_col99[45];
   data_col99[47] <= data_col99[46];
   data_col99[48] <= data_col99[47];
   data_col99[49] <= data_col99[48];
   data_col99[50] <= data_col99[49];
   data_col99[51] <= data_col99[50];
   data_col99[52] <= data_col99[51];
   data_col99[53] <= data_col99[52];
   data_col99[54] <= data_col99[53];
   data_col99[55] <= data_col99[54];
   data_col99[56] <= data_col99[55];
   data_col99[57] <= data_col99[56];
   data_col99[58] <= data_col99[57];
   data_col99[59] <= data_col99[58];
   data_col99[60] <= data_col99[59];
   data_col99[61] <= data_col99[60];
   data_col99[62] <= data_col99[61];
   data_col99[63] <= data_col99[62];
   data_col99[64] <= data_col99[63];
   data_col99[65] <= data_col99[64];
   data_col99[66] <= data_col99[65];
   data_col99[67] <= data_col99[66];
   data_col99[68] <= data_col99[67];
   data_col99[69] <= data_col99[68];
   data_col99[70] <= data_col99[69];
   data_col99[71] <= data_col99[70];
   data_col99[72] <= data_col99[71];
   data_col99[73] <= data_col99[72];
   data_col99[74] <= data_col99[73];
   data_col99[75] <= data_col99[74];
   data_col99[76] <= data_col99[75];
   data_col99[77] <= data_col99[76];
   data_col99[78] <= data_col99[77];
   data_col99[79] <= data_col99[78];
   data_col99[80] <= data_col99[79];
   data_col99[81] <= data_col99[80];
   data_col99[82] <= data_col99[81];
   data_col99[83] <= data_col99[82];
   data_col99[84] <= data_col99[83];
   data_col99[85] <= data_col99[84];
   data_col99[86] <= data_col99[85];
   data_col99[87] <= data_col99[86];
   data_col99[88] <= data_col99[87];
   data_col99[89] <= data_col99[88];
   data_col99[90] <= data_col99[89];
   data_col99[91] <= data_col99[90];
   data_col99[92] <= data_col99[91];
   data_col99[93] <= data_col99[92];
   data_col99[94] <= data_col99[93];
   data_col99[95] <= data_col99[94];
   data_col99[96] <= data_col99[95];
   data_col99[97] <= data_col99[96];
   data_col99[98] <= data_col99[97];
   data_col99[99] <= data_col99[98];

   data_col100[1] <= data[0];
   data_col100[2] <= data_col100[1];
   data_col100[3] <= data_col100[2];
   data_col100[4] <= data_col100[3];
   data_col100[5] <= data_col100[4];
   data_col100[6] <= data_col100[5];
   data_col100[7] <= data_col100[6];
   data_col100[8] <= data_col100[7];
   data_col100[9] <= data_col100[8];
   data_col100[10] <= data_col100[9];
   data_col100[11] <= data_col100[10];
   data_col100[12] <= data_col100[11];
   data_col100[13] <= data_col100[12];
   data_col100[14] <= data_col100[13];
   data_col100[15] <= data_col100[14];
   data_col100[16] <= data_col100[15];
   data_col100[17] <= data_col100[16];
   data_col100[18] <= data_col100[17];
   data_col100[19] <= data_col100[18];
   data_col100[20] <= data_col100[19];
   data_col100[21] <= data_col100[20];
   data_col100[22] <= data_col100[21];
   data_col100[23] <= data_col100[22];
   data_col100[24] <= data_col100[23];
   data_col100[25] <= data_col100[24];
   data_col100[26] <= data_col100[25];
   data_col100[27] <= data_col100[26];
   data_col100[28] <= data_col100[27];
   data_col100[29] <= data_col100[28];
   data_col100[30] <= data_col100[29];
   data_col100[31] <= data_col100[30];
   data_col100[32] <= data_col100[31];
   data_col100[33] <= data_col100[32];
   data_col100[34] <= data_col100[33];
   data_col100[35] <= data_col100[34];
   data_col100[36] <= data_col100[35];
   data_col100[37] <= data_col100[36];
   data_col100[38] <= data_col100[37];
   data_col100[39] <= data_col100[38];
   data_col100[40] <= data_col100[39];
   data_col100[41] <= data_col100[40];
   data_col100[42] <= data_col100[41];
   data_col100[43] <= data_col100[42];
   data_col100[44] <= data_col100[43];
   data_col100[45] <= data_col100[44];
   data_col100[46] <= data_col100[45];
   data_col100[47] <= data_col100[46];
   data_col100[48] <= data_col100[47];
   data_col100[49] <= data_col100[48];
   data_col100[50] <= data_col100[49];
   data_col100[51] <= data_col100[50];
   data_col100[52] <= data_col100[51];
   data_col100[53] <= data_col100[52];
   data_col100[54] <= data_col100[53];
   data_col100[55] <= data_col100[54];
   data_col100[56] <= data_col100[55];
   data_col100[57] <= data_col100[56];
   data_col100[58] <= data_col100[57];
   data_col100[59] <= data_col100[58];
   data_col100[60] <= data_col100[59];
   data_col100[61] <= data_col100[60];
   data_col100[62] <= data_col100[61];
   data_col100[63] <= data_col100[62];
   data_col100[64] <= data_col100[63];
   data_col100[65] <= data_col100[64];
   data_col100[66] <= data_col100[65];
   data_col100[67] <= data_col100[66];
   data_col100[68] <= data_col100[67];
   data_col100[69] <= data_col100[68];
   data_col100[70] <= data_col100[69];
   data_col100[71] <= data_col100[70];
   data_col100[72] <= data_col100[71];
   data_col100[73] <= data_col100[72];
   data_col100[74] <= data_col100[73];
   data_col100[75] <= data_col100[74];
   data_col100[76] <= data_col100[75];
   data_col100[77] <= data_col100[76];
   data_col100[78] <= data_col100[77];
   data_col100[79] <= data_col100[78];
   data_col100[80] <= data_col100[79];
   data_col100[81] <= data_col100[80];
   data_col100[82] <= data_col100[81];
   data_col100[83] <= data_col100[82];
   data_col100[84] <= data_col100[83];
   data_col100[85] <= data_col100[84];
   data_col100[86] <= data_col100[85];
   data_col100[87] <= data_col100[86];
   data_col100[88] <= data_col100[87];
   data_col100[89] <= data_col100[88];
   data_col100[90] <= data_col100[89];
   data_col100[91] <= data_col100[90];
   data_col100[92] <= data_col100[91];
   data_col100[93] <= data_col100[92];
   data_col100[94] <= data_col100[93];
   data_col100[95] <= data_col100[94];
   data_col100[96] <= data_col100[95];
   data_col100[97] <= data_col100[96];
   data_col100[98] <= data_col100[97];
   data_col100[99] <= data_col100[98];
   data_col100[100] <= data_col100[99];
 end

 wire [DAT_W-1:0] data_in;
 assign data_in = {data_col0, data_col1[1], data_col2[2], data_col3[3], data_col4[4], data_col5[5], data_col6[6], data_col7[7], data_col8[8], data_col9[9], data_col10[10], data_col11[11], data_col12[12], data_col13[13], data_col14[14], data_col15[15], data_col16[16], data_col17[17], data_col18[18], data_col19[19], data_col20[20], data_col21[21], data_col22[22], data_col23[23], data_col24[24], data_col25[25], data_col26[26], data_col27[27], data_col28[28], data_col29[29], data_col30[30], data_col31[31], data_col32[32], data_col33[33], data_col34[34], data_col35[35], data_col36[36], data_col37[37], data_col38[38], data_col39[39], data_col40[40], data_col41[41], data_col42[42], data_col43[43], data_col44[44], data_col45[45], data_col46[46], data_col47[47], data_col48[48], data_col49[49], data_col50[50], data_col51[51], data_col52[52], data_col53[53], data_col54[54], data_col55[55], data_col56[56], data_col57[57], data_col58[58], data_col59[59], data_col60[60], data_col61[61], data_col62[62], data_col63[63], data_col64[64], data_col65[65], data_col66[66], data_col67[67], data_col68[68], data_col69[69], data_col70[70], data_col71[71], data_col72[72], data_col73[73], data_col74[74], data_col75[75], data_col76[76], data_col77[77], data_col78[78], data_col79[79], data_col80[80], data_col81[81], data_col82[82], data_col83[83], data_col84[84], data_col85[85], data_col86[86], data_col87[87], data_col88[88], data_col89[89], data_col90[90], data_col91[91], data_col92[92], data_col93[93], data_col94[94], data_col95[95], data_col96[96], data_col97[97], data_col98[98], data_col99[99], data_col100[100]};

  /////////////////////////////////////
  // row 0
  // row 0, col 0

     wire start_in_0_0;
     wire start_out_0_0;

     wire [1:0] op_in_0_0;
     wire [1:0] op_out_0_0;

     wire r_0_0;

     wire data_in_0_0;
     wire data_out_0_0;

     wire pivot_in_0_0;
     wire pivot_out_0_0;

     assign data_in_0_0 = data_in[DAT_W-1];
     assign op_in_0_0 = mode & start ? 2'b01 : 2'b00;
     assign pivot_in_0_0 = 0;

     assign start_in_0_0 = start;

     processor_AB AB_0_0 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_0),
       .start_in   (start_in_0_0),
       .op_in      (op_in_0_0),
       .pivot_in   (pivot_in_0_0),
       .start_out  (start_out_0_0),
       .data_out   (data_out_0_0),
       .op_out     (op_out_0_0),
       .pivot_out  (pivot_out_0_0),
       .r          (r_0_0)
     );

  // row 0, col 1

     reg start_in_0_1;
     wire start_out_0_1;

     reg [1:0] op_in_0_1;
     wire [1:0] op_out_0_1;

     wire r_0_1;

     wire data_in_0_1;
     wire data_out_0_1;

     reg pivot_in_0_1;
     wire pivot_out_0_1;

     assign data_in_0_1 = data_in[DAT_W-2];

     always @(posedge clk) begin
        op_in_0_1 <= op_out_0_0;
        pivot_in_0_1 <= pivot_out_0_0;
        start_in_0_1 <= start_out_0_0;
     end
  
     processor_AB AB_0_1 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_1),
       .start_in   (start_in_0_1),
       .op_in      (op_in_0_1),
       .pivot_in   (pivot_in_0_1),
       .start_out  (start_out_0_1),
       .data_out   (data_out_0_1),
       .op_out     (op_out_0_1),
       .pivot_out  (pivot_out_0_1),
       .r          (r_0_1)
     );

  // row 0, col 2

     reg start_in_0_2;
     wire start_out_0_2;

     reg [1:0] op_in_0_2;
     wire [1:0] op_out_0_2;

     wire r_0_2;

     wire data_in_0_2;
     wire data_out_0_2;

     reg pivot_in_0_2;
     wire pivot_out_0_2;

     assign data_in_0_2 = data_in[DAT_W-3];

     always @(posedge clk) begin
        op_in_0_2 <= op_out_0_1;
        pivot_in_0_2 <= pivot_out_0_1;
        start_in_0_2 <= start_out_0_1;
     end
  
     processor_AB AB_0_2 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_2),
       .start_in   (start_in_0_2),
       .op_in      (op_in_0_2),
       .pivot_in   (pivot_in_0_2),
       .start_out  (start_out_0_2),
       .data_out   (data_out_0_2),
       .op_out     (op_out_0_2),
       .pivot_out  (pivot_out_0_2),
       .r          (r_0_2)
     );

  // row 0, col 3

     reg start_in_0_3;
     wire start_out_0_3;

     reg [1:0] op_in_0_3;
     wire [1:0] op_out_0_3;

     wire r_0_3;

     wire data_in_0_3;
     wire data_out_0_3;

     reg pivot_in_0_3;
     wire pivot_out_0_3;

     assign data_in_0_3 = data_in[DAT_W-4];

     always @(posedge clk) begin
        op_in_0_3 <= op_out_0_2;
        pivot_in_0_3 <= pivot_out_0_2;
        start_in_0_3 <= start_out_0_2;
     end
  
     processor_AB AB_0_3 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_3),
       .start_in   (start_in_0_3),
       .op_in      (op_in_0_3),
       .pivot_in   (pivot_in_0_3),
       .start_out  (start_out_0_3),
       .data_out   (data_out_0_3),
       .op_out     (op_out_0_3),
       .pivot_out  (pivot_out_0_3),
       .r          (r_0_3)
     );

  // row 0, col 4

     reg start_in_0_4;
     wire start_out_0_4;

     reg [1:0] op_in_0_4;
     wire [1:0] op_out_0_4;

     wire r_0_4;

     wire data_in_0_4;
     wire data_out_0_4;

     reg pivot_in_0_4;
     wire pivot_out_0_4;

     assign data_in_0_4 = data_in[DAT_W-5];

     always @(posedge clk) begin
        op_in_0_4 <= op_out_0_3;
        pivot_in_0_4 <= pivot_out_0_3;
        start_in_0_4 <= start_out_0_3;
     end
  
     processor_AB AB_0_4 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_4),
       .start_in   (start_in_0_4),
       .op_in      (op_in_0_4),
       .pivot_in   (pivot_in_0_4),
       .start_out  (start_out_0_4),
       .data_out   (data_out_0_4),
       .op_out     (op_out_0_4),
       .pivot_out  (pivot_out_0_4),
       .r          (r_0_4)
     );

  // row 0, col 5

     reg start_in_0_5;
     wire start_out_0_5;

     reg [1:0] op_in_0_5;
     wire [1:0] op_out_0_5;

     wire r_0_5;

     wire data_in_0_5;
     wire data_out_0_5;

     reg pivot_in_0_5;
     wire pivot_out_0_5;

     assign data_in_0_5 = data_in[DAT_W-6];

     always @(posedge clk) begin
        op_in_0_5 <= op_out_0_4;
        pivot_in_0_5 <= pivot_out_0_4;
        start_in_0_5 <= start_out_0_4;
     end
  
     processor_AB AB_0_5 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_5),
       .start_in   (start_in_0_5),
       .op_in      (op_in_0_5),
       .pivot_in   (pivot_in_0_5),
       .start_out  (start_out_0_5),
       .data_out   (data_out_0_5),
       .op_out     (op_out_0_5),
       .pivot_out  (pivot_out_0_5),
       .r          (r_0_5)
     );

  // row 0, col 6

     reg start_in_0_6;
     wire start_out_0_6;

     reg [1:0] op_in_0_6;
     wire [1:0] op_out_0_6;

     wire r_0_6;

     wire data_in_0_6;
     wire data_out_0_6;

     reg pivot_in_0_6;
     wire pivot_out_0_6;

     assign data_in_0_6 = data_in[DAT_W-7];

     always @(posedge clk) begin
        op_in_0_6 <= op_out_0_5;
        pivot_in_0_6 <= pivot_out_0_5;
        start_in_0_6 <= start_out_0_5;
     end
  
     processor_AB AB_0_6 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_6),
       .start_in   (start_in_0_6),
       .op_in      (op_in_0_6),
       .pivot_in   (pivot_in_0_6),
       .start_out  (start_out_0_6),
       .data_out   (data_out_0_6),
       .op_out     (op_out_0_6),
       .pivot_out  (pivot_out_0_6),
       .r          (r_0_6)
     );

  // row 0, col 7

     reg start_in_0_7;
     wire start_out_0_7;

     reg [1:0] op_in_0_7;
     wire [1:0] op_out_0_7;

     wire r_0_7;

     wire data_in_0_7;
     wire data_out_0_7;

     reg pivot_in_0_7;
     wire pivot_out_0_7;

     assign data_in_0_7 = data_in[DAT_W-8];

     always @(posedge clk) begin
        op_in_0_7 <= op_out_0_6;
        pivot_in_0_7 <= pivot_out_0_6;
        start_in_0_7 <= start_out_0_6;
     end
  
     processor_AB AB_0_7 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_7),
       .start_in   (start_in_0_7),
       .op_in      (op_in_0_7),
       .pivot_in   (pivot_in_0_7),
       .start_out  (start_out_0_7),
       .data_out   (data_out_0_7),
       .op_out     (op_out_0_7),
       .pivot_out  (pivot_out_0_7),
       .r          (r_0_7)
     );

  // row 0, col 8

     reg start_in_0_8;
     wire start_out_0_8;

     reg [1:0] op_in_0_8;
     wire [1:0] op_out_0_8;

     wire r_0_8;

     wire data_in_0_8;
     wire data_out_0_8;

     reg pivot_in_0_8;
     wire pivot_out_0_8;

     assign data_in_0_8 = data_in[DAT_W-9];

     always @(posedge clk) begin
        op_in_0_8 <= op_out_0_7;
        pivot_in_0_8 <= pivot_out_0_7;
        start_in_0_8 <= start_out_0_7;
     end
  
     processor_AB AB_0_8 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_8),
       .start_in   (start_in_0_8),
       .op_in      (op_in_0_8),
       .pivot_in   (pivot_in_0_8),
       .start_out  (start_out_0_8),
       .data_out   (data_out_0_8),
       .op_out     (op_out_0_8),
       .pivot_out  (pivot_out_0_8),
       .r          (r_0_8)
     );

  // row 0, col 9

     reg start_in_0_9;
     wire start_out_0_9;

     reg [1:0] op_in_0_9;
     wire [1:0] op_out_0_9;

     wire r_0_9;

     wire data_in_0_9;
     wire data_out_0_9;

     reg pivot_in_0_9;
     wire pivot_out_0_9;

     assign data_in_0_9 = data_in[DAT_W-10];

     always @(posedge clk) begin
        op_in_0_9 <= op_out_0_8;
        pivot_in_0_9 <= pivot_out_0_8;
        start_in_0_9 <= start_out_0_8;
     end
  
     processor_AB AB_0_9 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_9),
       .start_in   (start_in_0_9),
       .op_in      (op_in_0_9),
       .pivot_in   (pivot_in_0_9),
       .start_out  (start_out_0_9),
       .data_out   (data_out_0_9),
       .op_out     (op_out_0_9),
       .pivot_out  (pivot_out_0_9),
       .r          (r_0_9)
     );

  // row 0, col 10

     reg start_in_0_10;
     wire start_out_0_10;

     reg [1:0] op_in_0_10;
     wire [1:0] op_out_0_10;

     wire r_0_10;

     wire data_in_0_10;
     wire data_out_0_10;

     reg pivot_in_0_10;
     wire pivot_out_0_10;

     assign data_in_0_10 = data_in[DAT_W-11];

     always @(posedge clk) begin
        op_in_0_10 <= op_out_0_9;
        pivot_in_0_10 <= pivot_out_0_9;
        start_in_0_10 <= start_out_0_9;
     end
  
     processor_AB AB_0_10 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_10),
       .start_in   (start_in_0_10),
       .op_in      (op_in_0_10),
       .pivot_in   (pivot_in_0_10),
       .start_out  (start_out_0_10),
       .data_out   (data_out_0_10),
       .op_out     (op_out_0_10),
       .pivot_out  (pivot_out_0_10),
       .r          (r_0_10)
     );

  // row 0, col 11

     reg start_in_0_11;
     wire start_out_0_11;

     reg [1:0] op_in_0_11;
     wire [1:0] op_out_0_11;

     wire r_0_11;

     wire data_in_0_11;
     wire data_out_0_11;

     reg pivot_in_0_11;
     wire pivot_out_0_11;

     assign data_in_0_11 = data_in[DAT_W-12];

     always @(posedge clk) begin
        op_in_0_11 <= op_out_0_10;
        pivot_in_0_11 <= pivot_out_0_10;
        start_in_0_11 <= start_out_0_10;
     end
  
     processor_AB AB_0_11 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_11),
       .start_in   (start_in_0_11),
       .op_in      (op_in_0_11),
       .pivot_in   (pivot_in_0_11),
       .start_out  (start_out_0_11),
       .data_out   (data_out_0_11),
       .op_out     (op_out_0_11),
       .pivot_out  (pivot_out_0_11),
       .r          (r_0_11)
     );

  // row 0, col 12

     reg start_in_0_12;
     wire start_out_0_12;

     reg [1:0] op_in_0_12;
     wire [1:0] op_out_0_12;

     wire r_0_12;

     wire data_in_0_12;
     wire data_out_0_12;

     reg pivot_in_0_12;
     wire pivot_out_0_12;

     assign data_in_0_12 = data_in[DAT_W-13];

     always @(posedge clk) begin
        op_in_0_12 <= op_out_0_11;
        pivot_in_0_12 <= pivot_out_0_11;
        start_in_0_12 <= start_out_0_11;
     end
  
     processor_AB AB_0_12 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_12),
       .start_in   (start_in_0_12),
       .op_in      (op_in_0_12),
       .pivot_in   (pivot_in_0_12),
       .start_out  (start_out_0_12),
       .data_out   (data_out_0_12),
       .op_out     (op_out_0_12),
       .pivot_out  (pivot_out_0_12),
       .r          (r_0_12)
     );

  // row 0, col 13

     reg start_in_0_13;
     wire start_out_0_13;

     reg [1:0] op_in_0_13;
     wire [1:0] op_out_0_13;

     wire r_0_13;

     wire data_in_0_13;
     wire data_out_0_13;

     reg pivot_in_0_13;
     wire pivot_out_0_13;

     assign data_in_0_13 = data_in[DAT_W-14];

     always @(posedge clk) begin
        op_in_0_13 <= op_out_0_12;
        pivot_in_0_13 <= pivot_out_0_12;
        start_in_0_13 <= start_out_0_12;
     end
  
     processor_AB AB_0_13 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_13),
       .start_in   (start_in_0_13),
       .op_in      (op_in_0_13),
       .pivot_in   (pivot_in_0_13),
       .start_out  (start_out_0_13),
       .data_out   (data_out_0_13),
       .op_out     (op_out_0_13),
       .pivot_out  (pivot_out_0_13),
       .r          (r_0_13)
     );

  // row 0, col 14

     reg start_in_0_14;
     wire start_out_0_14;

     reg [1:0] op_in_0_14;
     wire [1:0] op_out_0_14;

     wire r_0_14;

     wire data_in_0_14;
     wire data_out_0_14;

     reg pivot_in_0_14;
     wire pivot_out_0_14;

     assign data_in_0_14 = data_in[DAT_W-15];

     always @(posedge clk) begin
        op_in_0_14 <= op_out_0_13;
        pivot_in_0_14 <= pivot_out_0_13;
        start_in_0_14 <= start_out_0_13;
     end
  
     processor_AB AB_0_14 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_14),
       .start_in   (start_in_0_14),
       .op_in      (op_in_0_14),
       .pivot_in   (pivot_in_0_14),
       .start_out  (start_out_0_14),
       .data_out   (data_out_0_14),
       .op_out     (op_out_0_14),
       .pivot_out  (pivot_out_0_14),
       .r          (r_0_14)
     );

  // row 0, col 15

     reg start_in_0_15;
     wire start_out_0_15;

     reg [1:0] op_in_0_15;
     wire [1:0] op_out_0_15;

     wire r_0_15;

     wire data_in_0_15;
     wire data_out_0_15;

     reg pivot_in_0_15;
     wire pivot_out_0_15;

     assign data_in_0_15 = data_in[DAT_W-16];

     always @(posedge clk) begin
        op_in_0_15 <= op_out_0_14;
        pivot_in_0_15 <= pivot_out_0_14;
        start_in_0_15 <= start_out_0_14;
     end
  
     processor_AB AB_0_15 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_15),
       .start_in   (start_in_0_15),
       .op_in      (op_in_0_15),
       .pivot_in   (pivot_in_0_15),
       .start_out  (start_out_0_15),
       .data_out   (data_out_0_15),
       .op_out     (op_out_0_15),
       .pivot_out  (pivot_out_0_15),
       .r          (r_0_15)
     );

  // row 0, col 16

     reg start_in_0_16;
     wire start_out_0_16;

     reg [1:0] op_in_0_16;
     wire [1:0] op_out_0_16;

     wire r_0_16;

     wire data_in_0_16;
     wire data_out_0_16;

     reg pivot_in_0_16;
     wire pivot_out_0_16;

     assign data_in_0_16 = data_in[DAT_W-17];

     always @(posedge clk) begin
        op_in_0_16 <= op_out_0_15;
        pivot_in_0_16 <= pivot_out_0_15;
        start_in_0_16 <= start_out_0_15;
     end
  
     processor_AB AB_0_16 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_16),
       .start_in   (start_in_0_16),
       .op_in      (op_in_0_16),
       .pivot_in   (pivot_in_0_16),
       .start_out  (start_out_0_16),
       .data_out   (data_out_0_16),
       .op_out     (op_out_0_16),
       .pivot_out  (pivot_out_0_16),
       .r          (r_0_16)
     );

  // row 0, col 17

     reg start_in_0_17;
     wire start_out_0_17;

     reg [1:0] op_in_0_17;
     wire [1:0] op_out_0_17;

     wire r_0_17;

     wire data_in_0_17;
     wire data_out_0_17;

     reg pivot_in_0_17;
     wire pivot_out_0_17;

     assign data_in_0_17 = data_in[DAT_W-18];

     always @(posedge clk) begin
        op_in_0_17 <= op_out_0_16;
        pivot_in_0_17 <= pivot_out_0_16;
        start_in_0_17 <= start_out_0_16;
     end
  
     processor_AB AB_0_17 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_17),
       .start_in   (start_in_0_17),
       .op_in      (op_in_0_17),
       .pivot_in   (pivot_in_0_17),
       .start_out  (start_out_0_17),
       .data_out   (data_out_0_17),
       .op_out     (op_out_0_17),
       .pivot_out  (pivot_out_0_17),
       .r          (r_0_17)
     );

  // row 0, col 18

     reg start_in_0_18;
     wire start_out_0_18;

     reg [1:0] op_in_0_18;
     wire [1:0] op_out_0_18;

     wire r_0_18;

     wire data_in_0_18;
     wire data_out_0_18;

     reg pivot_in_0_18;
     wire pivot_out_0_18;

     assign data_in_0_18 = data_in[DAT_W-19];

     always @(posedge clk) begin
        op_in_0_18 <= op_out_0_17;
        pivot_in_0_18 <= pivot_out_0_17;
        start_in_0_18 <= start_out_0_17;
     end
  
     processor_AB AB_0_18 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_18),
       .start_in   (start_in_0_18),
       .op_in      (op_in_0_18),
       .pivot_in   (pivot_in_0_18),
       .start_out  (start_out_0_18),
       .data_out   (data_out_0_18),
       .op_out     (op_out_0_18),
       .pivot_out  (pivot_out_0_18),
       .r          (r_0_18)
     );

  // row 0, col 19

     reg start_in_0_19;
     wire start_out_0_19;

     reg [1:0] op_in_0_19;
     wire [1:0] op_out_0_19;

     wire r_0_19;

     wire data_in_0_19;
     wire data_out_0_19;

     reg pivot_in_0_19;
     wire pivot_out_0_19;

     assign data_in_0_19 = data_in[DAT_W-20];

     always @(posedge clk) begin
        op_in_0_19 <= op_out_0_18;
        pivot_in_0_19 <= pivot_out_0_18;
        start_in_0_19 <= start_out_0_18;
     end
  
     processor_AB AB_0_19 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_19),
       .start_in   (start_in_0_19),
       .op_in      (op_in_0_19),
       .pivot_in   (pivot_in_0_19),
       .start_out  (start_out_0_19),
       .data_out   (data_out_0_19),
       .op_out     (op_out_0_19),
       .pivot_out  (pivot_out_0_19),
       .r          (r_0_19)
     );

  // row 0, col 20

     reg start_in_0_20;
     wire start_out_0_20;

     reg [1:0] op_in_0_20;
     wire [1:0] op_out_0_20;

     wire r_0_20;

     wire data_in_0_20;
     wire data_out_0_20;

     reg pivot_in_0_20;
     wire pivot_out_0_20;

     assign data_in_0_20 = data_in[DAT_W-21];

     always @(posedge clk) begin
        op_in_0_20 <= op_out_0_19;
        pivot_in_0_20 <= pivot_out_0_19;
        start_in_0_20 <= start_out_0_19;
     end
  
     processor_AB AB_0_20 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_20),
       .start_in   (start_in_0_20),
       .op_in      (op_in_0_20),
       .pivot_in   (pivot_in_0_20),
       .start_out  (start_out_0_20),
       .data_out   (data_out_0_20),
       .op_out     (op_out_0_20),
       .pivot_out  (pivot_out_0_20),
       .r          (r_0_20)
     );

  // row 0, col 21

     reg start_in_0_21;
     wire start_out_0_21;

     reg [1:0] op_in_0_21;
     wire [1:0] op_out_0_21;

     wire r_0_21;

     wire data_in_0_21;
     wire data_out_0_21;

     reg pivot_in_0_21;
     wire pivot_out_0_21;

     assign data_in_0_21 = data_in[DAT_W-22];

     always @(posedge clk) begin
        op_in_0_21 <= op_out_0_20;
        pivot_in_0_21 <= pivot_out_0_20;
        start_in_0_21 <= start_out_0_20;
     end
  
     processor_AB AB_0_21 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_21),
       .start_in   (start_in_0_21),
       .op_in      (op_in_0_21),
       .pivot_in   (pivot_in_0_21),
       .start_out  (start_out_0_21),
       .data_out   (data_out_0_21),
       .op_out     (op_out_0_21),
       .pivot_out  (pivot_out_0_21),
       .r          (r_0_21)
     );

  // row 0, col 22

     reg start_in_0_22;
     wire start_out_0_22;

     reg [1:0] op_in_0_22;
     wire [1:0] op_out_0_22;

     wire r_0_22;

     wire data_in_0_22;
     wire data_out_0_22;

     reg pivot_in_0_22;
     wire pivot_out_0_22;

     assign data_in_0_22 = data_in[DAT_W-23];

     always @(posedge clk) begin
        op_in_0_22 <= op_out_0_21;
        pivot_in_0_22 <= pivot_out_0_21;
        start_in_0_22 <= start_out_0_21;
     end
  
     processor_AB AB_0_22 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_22),
       .start_in   (start_in_0_22),
       .op_in      (op_in_0_22),
       .pivot_in   (pivot_in_0_22),
       .start_out  (start_out_0_22),
       .data_out   (data_out_0_22),
       .op_out     (op_out_0_22),
       .pivot_out  (pivot_out_0_22),
       .r          (r_0_22)
     );

  // row 0, col 23

     reg start_in_0_23;
     wire start_out_0_23;

     reg [1:0] op_in_0_23;
     wire [1:0] op_out_0_23;

     wire r_0_23;

     wire data_in_0_23;
     wire data_out_0_23;

     reg pivot_in_0_23;
     wire pivot_out_0_23;

     assign data_in_0_23 = data_in[DAT_W-24];

     always @(posedge clk) begin
        op_in_0_23 <= op_out_0_22;
        pivot_in_0_23 <= pivot_out_0_22;
        start_in_0_23 <= start_out_0_22;
     end
  
     processor_AB AB_0_23 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_23),
       .start_in   (start_in_0_23),
       .op_in      (op_in_0_23),
       .pivot_in   (pivot_in_0_23),
       .start_out  (start_out_0_23),
       .data_out   (data_out_0_23),
       .op_out     (op_out_0_23),
       .pivot_out  (pivot_out_0_23),
       .r          (r_0_23)
     );

  // row 0, col 24

     reg start_in_0_24;
     wire start_out_0_24;

     reg [1:0] op_in_0_24;
     wire [1:0] op_out_0_24;

     wire r_0_24;

     wire data_in_0_24;
     wire data_out_0_24;

     reg pivot_in_0_24;
     wire pivot_out_0_24;

     assign data_in_0_24 = data_in[DAT_W-25];

     always @(posedge clk) begin
        op_in_0_24 <= op_out_0_23;
        pivot_in_0_24 <= pivot_out_0_23;
        start_in_0_24 <= start_out_0_23;
     end
  
     processor_AB AB_0_24 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_24),
       .start_in   (start_in_0_24),
       .op_in      (op_in_0_24),
       .pivot_in   (pivot_in_0_24),
       .start_out  (start_out_0_24),
       .data_out   (data_out_0_24),
       .op_out     (op_out_0_24),
       .pivot_out  (pivot_out_0_24),
       .r          (r_0_24)
     );

  // row 0, col 25

     reg start_in_0_25;
     wire start_out_0_25;

     reg [1:0] op_in_0_25;
     wire [1:0] op_out_0_25;

     wire r_0_25;

     wire data_in_0_25;
     wire data_out_0_25;

     reg pivot_in_0_25;
     wire pivot_out_0_25;

     assign data_in_0_25 = data_in[DAT_W-26];

     always @(posedge clk) begin
        op_in_0_25 <= op_out_0_24;
        pivot_in_0_25 <= pivot_out_0_24;
        start_in_0_25 <= start_out_0_24;
     end
  
     processor_AB AB_0_25 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_25),
       .start_in   (start_in_0_25),
       .op_in      (op_in_0_25),
       .pivot_in   (pivot_in_0_25),
       .start_out  (start_out_0_25),
       .data_out   (data_out_0_25),
       .op_out     (op_out_0_25),
       .pivot_out  (pivot_out_0_25),
       .r          (r_0_25)
     );

  // row 0, col 26

     reg start_in_0_26;
     wire start_out_0_26;

     reg [1:0] op_in_0_26;
     wire [1:0] op_out_0_26;

     wire r_0_26;

     wire data_in_0_26;
     wire data_out_0_26;

     reg pivot_in_0_26;
     wire pivot_out_0_26;

     assign data_in_0_26 = data_in[DAT_W-27];

     always @(posedge clk) begin
        op_in_0_26 <= op_out_0_25;
        pivot_in_0_26 <= pivot_out_0_25;
        start_in_0_26 <= start_out_0_25;
     end
  
     processor_AB AB_0_26 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_26),
       .start_in   (start_in_0_26),
       .op_in      (op_in_0_26),
       .pivot_in   (pivot_in_0_26),
       .start_out  (start_out_0_26),
       .data_out   (data_out_0_26),
       .op_out     (op_out_0_26),
       .pivot_out  (pivot_out_0_26),
       .r          (r_0_26)
     );

  // row 0, col 27

     reg start_in_0_27;
     wire start_out_0_27;

     reg [1:0] op_in_0_27;
     wire [1:0] op_out_0_27;

     wire r_0_27;

     wire data_in_0_27;
     wire data_out_0_27;

     reg pivot_in_0_27;
     wire pivot_out_0_27;

     assign data_in_0_27 = data_in[DAT_W-28];

     always @(posedge clk) begin
        op_in_0_27 <= op_out_0_26;
        pivot_in_0_27 <= pivot_out_0_26;
        start_in_0_27 <= start_out_0_26;
     end
  
     processor_AB AB_0_27 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_27),
       .start_in   (start_in_0_27),
       .op_in      (op_in_0_27),
       .pivot_in   (pivot_in_0_27),
       .start_out  (start_out_0_27),
       .data_out   (data_out_0_27),
       .op_out     (op_out_0_27),
       .pivot_out  (pivot_out_0_27),
       .r          (r_0_27)
     );

  // row 0, col 28

     reg start_in_0_28;
     wire start_out_0_28;

     reg [1:0] op_in_0_28;
     wire [1:0] op_out_0_28;

     wire r_0_28;

     wire data_in_0_28;
     wire data_out_0_28;

     reg pivot_in_0_28;
     wire pivot_out_0_28;

     assign data_in_0_28 = data_in[DAT_W-29];

     always @(posedge clk) begin
        op_in_0_28 <= op_out_0_27;
        pivot_in_0_28 <= pivot_out_0_27;
        start_in_0_28 <= start_out_0_27;
     end
  
     processor_AB AB_0_28 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_28),
       .start_in   (start_in_0_28),
       .op_in      (op_in_0_28),
       .pivot_in   (pivot_in_0_28),
       .start_out  (start_out_0_28),
       .data_out   (data_out_0_28),
       .op_out     (op_out_0_28),
       .pivot_out  (pivot_out_0_28),
       .r          (r_0_28)
     );

  // row 0, col 29

     reg start_in_0_29;
     wire start_out_0_29;

     reg [1:0] op_in_0_29;
     wire [1:0] op_out_0_29;

     wire r_0_29;

     wire data_in_0_29;
     wire data_out_0_29;

     reg pivot_in_0_29;
     wire pivot_out_0_29;

     assign data_in_0_29 = data_in[DAT_W-30];

     always @(posedge clk) begin
        op_in_0_29 <= op_out_0_28;
        pivot_in_0_29 <= pivot_out_0_28;
        start_in_0_29 <= start_out_0_28;
     end
  
     processor_AB AB_0_29 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_29),
       .start_in   (start_in_0_29),
       .op_in      (op_in_0_29),
       .pivot_in   (pivot_in_0_29),
       .start_out  (start_out_0_29),
       .data_out   (data_out_0_29),
       .op_out     (op_out_0_29),
       .pivot_out  (pivot_out_0_29),
       .r          (r_0_29)
     );

  // row 0, col 30

     reg start_in_0_30;
     wire start_out_0_30;

     reg [1:0] op_in_0_30;
     wire [1:0] op_out_0_30;

     wire r_0_30;

     wire data_in_0_30;
     wire data_out_0_30;

     reg pivot_in_0_30;
     wire pivot_out_0_30;

     assign data_in_0_30 = data_in[DAT_W-31];

     always @(posedge clk) begin
        op_in_0_30 <= op_out_0_29;
        pivot_in_0_30 <= pivot_out_0_29;
        start_in_0_30 <= start_out_0_29;
     end
  
     processor_AB AB_0_30 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_30),
       .start_in   (start_in_0_30),
       .op_in      (op_in_0_30),
       .pivot_in   (pivot_in_0_30),
       .start_out  (start_out_0_30),
       .data_out   (data_out_0_30),
       .op_out     (op_out_0_30),
       .pivot_out  (pivot_out_0_30),
       .r          (r_0_30)
     );

  // row 0, col 31

     reg start_in_0_31;
     wire start_out_0_31;

     reg [1:0] op_in_0_31;
     wire [1:0] op_out_0_31;

     wire r_0_31;

     wire data_in_0_31;
     wire data_out_0_31;

     reg pivot_in_0_31;
     wire pivot_out_0_31;

     assign data_in_0_31 = data_in[DAT_W-32];

     always @(posedge clk) begin
        op_in_0_31 <= op_out_0_30;
        pivot_in_0_31 <= pivot_out_0_30;
        start_in_0_31 <= start_out_0_30;
     end
  
     processor_AB AB_0_31 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_31),
       .start_in   (start_in_0_31),
       .op_in      (op_in_0_31),
       .pivot_in   (pivot_in_0_31),
       .start_out  (start_out_0_31),
       .data_out   (data_out_0_31),
       .op_out     (op_out_0_31),
       .pivot_out  (pivot_out_0_31),
       .r          (r_0_31)
     );

  // row 0, col 32

     reg start_in_0_32;
     wire start_out_0_32;

     reg [1:0] op_in_0_32;
     wire [1:0] op_out_0_32;

     wire r_0_32;

     wire data_in_0_32;
     wire data_out_0_32;

     reg pivot_in_0_32;
     wire pivot_out_0_32;

     assign data_in_0_32 = data_in[DAT_W-33];

     always @(posedge clk) begin
        op_in_0_32 <= op_out_0_31;
        pivot_in_0_32 <= pivot_out_0_31;
        start_in_0_32 <= start_out_0_31;
     end
  
     processor_AB AB_0_32 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_32),
       .start_in   (start_in_0_32),
       .op_in      (op_in_0_32),
       .pivot_in   (pivot_in_0_32),
       .start_out  (start_out_0_32),
       .data_out   (data_out_0_32),
       .op_out     (op_out_0_32),
       .pivot_out  (pivot_out_0_32),
       .r          (r_0_32)
     );

  // row 0, col 33

     reg start_in_0_33;
     wire start_out_0_33;

     reg [1:0] op_in_0_33;
     wire [1:0] op_out_0_33;

     wire r_0_33;

     wire data_in_0_33;
     wire data_out_0_33;

     reg pivot_in_0_33;
     wire pivot_out_0_33;

     assign data_in_0_33 = data_in[DAT_W-34];

     always @(posedge clk) begin
        op_in_0_33 <= op_out_0_32;
        pivot_in_0_33 <= pivot_out_0_32;
        start_in_0_33 <= start_out_0_32;
     end
  
     processor_AB AB_0_33 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_33),
       .start_in   (start_in_0_33),
       .op_in      (op_in_0_33),
       .pivot_in   (pivot_in_0_33),
       .start_out  (start_out_0_33),
       .data_out   (data_out_0_33),
       .op_out     (op_out_0_33),
       .pivot_out  (pivot_out_0_33),
       .r          (r_0_33)
     );

  // row 0, col 34

     reg start_in_0_34;
     wire start_out_0_34;

     reg [1:0] op_in_0_34;
     wire [1:0] op_out_0_34;

     wire r_0_34;

     wire data_in_0_34;
     wire data_out_0_34;

     reg pivot_in_0_34;
     wire pivot_out_0_34;

     assign data_in_0_34 = data_in[DAT_W-35];

     always @(posedge clk) begin
        op_in_0_34 <= op_out_0_33;
        pivot_in_0_34 <= pivot_out_0_33;
        start_in_0_34 <= start_out_0_33;
     end
  
     processor_AB AB_0_34 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_34),
       .start_in   (start_in_0_34),
       .op_in      (op_in_0_34),
       .pivot_in   (pivot_in_0_34),
       .start_out  (start_out_0_34),
       .data_out   (data_out_0_34),
       .op_out     (op_out_0_34),
       .pivot_out  (pivot_out_0_34),
       .r          (r_0_34)
     );

  // row 0, col 35

     reg start_in_0_35;
     wire start_out_0_35;

     reg [1:0] op_in_0_35;
     wire [1:0] op_out_0_35;

     wire r_0_35;

     wire data_in_0_35;
     wire data_out_0_35;

     reg pivot_in_0_35;
     wire pivot_out_0_35;

     assign data_in_0_35 = data_in[DAT_W-36];

     always @(posedge clk) begin
        op_in_0_35 <= op_out_0_34;
        pivot_in_0_35 <= pivot_out_0_34;
        start_in_0_35 <= start_out_0_34;
     end
  
     processor_AB AB_0_35 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_35),
       .start_in   (start_in_0_35),
       .op_in      (op_in_0_35),
       .pivot_in   (pivot_in_0_35),
       .start_out  (start_out_0_35),
       .data_out   (data_out_0_35),
       .op_out     (op_out_0_35),
       .pivot_out  (pivot_out_0_35),
       .r          (r_0_35)
     );

  // row 0, col 36

     reg start_in_0_36;
     wire start_out_0_36;

     reg [1:0] op_in_0_36;
     wire [1:0] op_out_0_36;

     wire r_0_36;

     wire data_in_0_36;
     wire data_out_0_36;

     reg pivot_in_0_36;
     wire pivot_out_0_36;

     assign data_in_0_36 = data_in[DAT_W-37];

     always @(posedge clk) begin
        op_in_0_36 <= op_out_0_35;
        pivot_in_0_36 <= pivot_out_0_35;
        start_in_0_36 <= start_out_0_35;
     end
  
     processor_AB AB_0_36 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_36),
       .start_in   (start_in_0_36),
       .op_in      (op_in_0_36),
       .pivot_in   (pivot_in_0_36),
       .start_out  (start_out_0_36),
       .data_out   (data_out_0_36),
       .op_out     (op_out_0_36),
       .pivot_out  (pivot_out_0_36),
       .r          (r_0_36)
     );

  // row 0, col 37

     reg start_in_0_37;
     wire start_out_0_37;

     reg [1:0] op_in_0_37;
     wire [1:0] op_out_0_37;

     wire r_0_37;

     wire data_in_0_37;
     wire data_out_0_37;

     reg pivot_in_0_37;
     wire pivot_out_0_37;

     assign data_in_0_37 = data_in[DAT_W-38];

     always @(posedge clk) begin
        op_in_0_37 <= op_out_0_36;
        pivot_in_0_37 <= pivot_out_0_36;
        start_in_0_37 <= start_out_0_36;
     end
  
     processor_AB AB_0_37 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_37),
       .start_in   (start_in_0_37),
       .op_in      (op_in_0_37),
       .pivot_in   (pivot_in_0_37),
       .start_out  (start_out_0_37),
       .data_out   (data_out_0_37),
       .op_out     (op_out_0_37),
       .pivot_out  (pivot_out_0_37),
       .r          (r_0_37)
     );

  // row 0, col 38

     reg start_in_0_38;
     wire start_out_0_38;

     reg [1:0] op_in_0_38;
     wire [1:0] op_out_0_38;

     wire r_0_38;

     wire data_in_0_38;
     wire data_out_0_38;

     reg pivot_in_0_38;
     wire pivot_out_0_38;

     assign data_in_0_38 = data_in[DAT_W-39];

     always @(posedge clk) begin
        op_in_0_38 <= op_out_0_37;
        pivot_in_0_38 <= pivot_out_0_37;
        start_in_0_38 <= start_out_0_37;
     end
  
     processor_AB AB_0_38 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_38),
       .start_in   (start_in_0_38),
       .op_in      (op_in_0_38),
       .pivot_in   (pivot_in_0_38),
       .start_out  (start_out_0_38),
       .data_out   (data_out_0_38),
       .op_out     (op_out_0_38),
       .pivot_out  (pivot_out_0_38),
       .r          (r_0_38)
     );

  // row 0, col 39

     reg start_in_0_39;
     wire start_out_0_39;

     reg [1:0] op_in_0_39;
     wire [1:0] op_out_0_39;

     wire r_0_39;

     wire data_in_0_39;
     wire data_out_0_39;

     reg pivot_in_0_39;
     wire pivot_out_0_39;

     assign data_in_0_39 = data_in[DAT_W-40];

     always @(posedge clk) begin
        op_in_0_39 <= op_out_0_38;
        pivot_in_0_39 <= pivot_out_0_38;
        start_in_0_39 <= start_out_0_38;
     end
  
     processor_AB AB_0_39 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_39),
       .start_in   (start_in_0_39),
       .op_in      (op_in_0_39),
       .pivot_in   (pivot_in_0_39),
       .start_out  (start_out_0_39),
       .data_out   (data_out_0_39),
       .op_out     (op_out_0_39),
       .pivot_out  (pivot_out_0_39),
       .r          (r_0_39)
     );

  // row 0, col 40

     reg start_in_0_40;
     wire start_out_0_40;

     reg [1:0] op_in_0_40;
     wire [1:0] op_out_0_40;

     wire r_0_40;

     wire data_in_0_40;
     wire data_out_0_40;

     reg pivot_in_0_40;
     wire pivot_out_0_40;

     assign data_in_0_40 = data_in[DAT_W-41];

     always @(posedge clk) begin
        op_in_0_40 <= op_out_0_39;
        pivot_in_0_40 <= pivot_out_0_39;
        start_in_0_40 <= start_out_0_39;
     end
  
     processor_AB AB_0_40 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_40),
       .start_in   (start_in_0_40),
       .op_in      (op_in_0_40),
       .pivot_in   (pivot_in_0_40),
       .start_out  (start_out_0_40),
       .data_out   (data_out_0_40),
       .op_out     (op_out_0_40),
       .pivot_out  (pivot_out_0_40),
       .r          (r_0_40)
     );

  // row 0, col 41

     reg start_in_0_41;
     wire start_out_0_41;

     reg [1:0] op_in_0_41;
     wire [1:0] op_out_0_41;

     wire r_0_41;

     wire data_in_0_41;
     wire data_out_0_41;

     reg pivot_in_0_41;
     wire pivot_out_0_41;

     assign data_in_0_41 = data_in[DAT_W-42];

     always @(posedge clk) begin
        op_in_0_41 <= op_out_0_40;
        pivot_in_0_41 <= pivot_out_0_40;
        start_in_0_41 <= start_out_0_40;
     end
  
     processor_AB AB_0_41 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_41),
       .start_in   (start_in_0_41),
       .op_in      (op_in_0_41),
       .pivot_in   (pivot_in_0_41),
       .start_out  (start_out_0_41),
       .data_out   (data_out_0_41),
       .op_out     (op_out_0_41),
       .pivot_out  (pivot_out_0_41),
       .r          (r_0_41)
     );

  // row 0, col 42

     reg start_in_0_42;
     wire start_out_0_42;

     reg [1:0] op_in_0_42;
     wire [1:0] op_out_0_42;

     wire r_0_42;

     wire data_in_0_42;
     wire data_out_0_42;

     reg pivot_in_0_42;
     wire pivot_out_0_42;

     assign data_in_0_42 = data_in[DAT_W-43];

     always @(posedge clk) begin
        op_in_0_42 <= op_out_0_41;
        pivot_in_0_42 <= pivot_out_0_41;
        start_in_0_42 <= start_out_0_41;
     end
  
     processor_AB AB_0_42 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_42),
       .start_in   (start_in_0_42),
       .op_in      (op_in_0_42),
       .pivot_in   (pivot_in_0_42),
       .start_out  (start_out_0_42),
       .data_out   (data_out_0_42),
       .op_out     (op_out_0_42),
       .pivot_out  (pivot_out_0_42),
       .r          (r_0_42)
     );

  // row 0, col 43

     reg start_in_0_43;
     wire start_out_0_43;

     reg [1:0] op_in_0_43;
     wire [1:0] op_out_0_43;

     wire r_0_43;

     wire data_in_0_43;
     wire data_out_0_43;

     reg pivot_in_0_43;
     wire pivot_out_0_43;

     assign data_in_0_43 = data_in[DAT_W-44];

     always @(posedge clk) begin
        op_in_0_43 <= op_out_0_42;
        pivot_in_0_43 <= pivot_out_0_42;
        start_in_0_43 <= start_out_0_42;
     end
  
     processor_AB AB_0_43 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_43),
       .start_in   (start_in_0_43),
       .op_in      (op_in_0_43),
       .pivot_in   (pivot_in_0_43),
       .start_out  (start_out_0_43),
       .data_out   (data_out_0_43),
       .op_out     (op_out_0_43),
       .pivot_out  (pivot_out_0_43),
       .r          (r_0_43)
     );

  // row 0, col 44

     reg start_in_0_44;
     wire start_out_0_44;

     reg [1:0] op_in_0_44;
     wire [1:0] op_out_0_44;

     wire r_0_44;

     wire data_in_0_44;
     wire data_out_0_44;

     reg pivot_in_0_44;
     wire pivot_out_0_44;

     assign data_in_0_44 = data_in[DAT_W-45];

     always @(posedge clk) begin
        op_in_0_44 <= op_out_0_43;
        pivot_in_0_44 <= pivot_out_0_43;
        start_in_0_44 <= start_out_0_43;
     end
  
     processor_AB AB_0_44 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_44),
       .start_in   (start_in_0_44),
       .op_in      (op_in_0_44),
       .pivot_in   (pivot_in_0_44),
       .start_out  (start_out_0_44),
       .data_out   (data_out_0_44),
       .op_out     (op_out_0_44),
       .pivot_out  (pivot_out_0_44),
       .r          (r_0_44)
     );

  // row 0, col 45

     reg start_in_0_45;
     wire start_out_0_45;

     reg [1:0] op_in_0_45;
     wire [1:0] op_out_0_45;

     wire r_0_45;

     wire data_in_0_45;
     wire data_out_0_45;

     reg pivot_in_0_45;
     wire pivot_out_0_45;

     assign data_in_0_45 = data_in[DAT_W-46];

     always @(posedge clk) begin
        op_in_0_45 <= op_out_0_44;
        pivot_in_0_45 <= pivot_out_0_44;
        start_in_0_45 <= start_out_0_44;
     end
  
     processor_AB AB_0_45 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_45),
       .start_in   (start_in_0_45),
       .op_in      (op_in_0_45),
       .pivot_in   (pivot_in_0_45),
       .start_out  (start_out_0_45),
       .data_out   (data_out_0_45),
       .op_out     (op_out_0_45),
       .pivot_out  (pivot_out_0_45),
       .r          (r_0_45)
     );

  // row 0, col 46

     reg start_in_0_46;
     wire start_out_0_46;

     reg [1:0] op_in_0_46;
     wire [1:0] op_out_0_46;

     wire r_0_46;

     wire data_in_0_46;
     wire data_out_0_46;

     reg pivot_in_0_46;
     wire pivot_out_0_46;

     assign data_in_0_46 = data_in[DAT_W-47];

     always @(posedge clk) begin
        op_in_0_46 <= op_out_0_45;
        pivot_in_0_46 <= pivot_out_0_45;
        start_in_0_46 <= start_out_0_45;
     end
  
     processor_AB AB_0_46 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_46),
       .start_in   (start_in_0_46),
       .op_in      (op_in_0_46),
       .pivot_in   (pivot_in_0_46),
       .start_out  (start_out_0_46),
       .data_out   (data_out_0_46),
       .op_out     (op_out_0_46),
       .pivot_out  (pivot_out_0_46),
       .r          (r_0_46)
     );

  // row 0, col 47

     reg start_in_0_47;
     wire start_out_0_47;

     reg [1:0] op_in_0_47;
     wire [1:0] op_out_0_47;

     wire r_0_47;

     wire data_in_0_47;
     wire data_out_0_47;

     reg pivot_in_0_47;
     wire pivot_out_0_47;

     assign data_in_0_47 = data_in[DAT_W-48];

     always @(posedge clk) begin
        op_in_0_47 <= op_out_0_46;
        pivot_in_0_47 <= pivot_out_0_46;
        start_in_0_47 <= start_out_0_46;
     end
  
     processor_AB AB_0_47 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_47),
       .start_in   (start_in_0_47),
       .op_in      (op_in_0_47),
       .pivot_in   (pivot_in_0_47),
       .start_out  (start_out_0_47),
       .data_out   (data_out_0_47),
       .op_out     (op_out_0_47),
       .pivot_out  (pivot_out_0_47),
       .r          (r_0_47)
     );

  // row 0, col 48

     reg start_in_0_48;
     wire start_out_0_48;

     reg [1:0] op_in_0_48;
     wire [1:0] op_out_0_48;

     wire r_0_48;

     wire data_in_0_48;
     wire data_out_0_48;

     reg pivot_in_0_48;
     wire pivot_out_0_48;

     assign data_in_0_48 = data_in[DAT_W-49];

     always @(posedge clk) begin
        op_in_0_48 <= op_out_0_47;
        pivot_in_0_48 <= pivot_out_0_47;
        start_in_0_48 <= start_out_0_47;
     end
  
     processor_AB AB_0_48 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_48),
       .start_in   (start_in_0_48),
       .op_in      (op_in_0_48),
       .pivot_in   (pivot_in_0_48),
       .start_out  (start_out_0_48),
       .data_out   (data_out_0_48),
       .op_out     (op_out_0_48),
       .pivot_out  (pivot_out_0_48),
       .r          (r_0_48)
     );

  // row 0, col 49

     reg start_in_0_49;
     wire start_out_0_49;

     reg [1:0] op_in_0_49;
     wire [1:0] op_out_0_49;

     wire r_0_49;

     wire data_in_0_49;
     wire data_out_0_49;

     reg pivot_in_0_49;
     wire pivot_out_0_49;

     assign data_in_0_49 = data_in[DAT_W-50];

     always @(posedge clk) begin
        op_in_0_49 <= op_out_0_48;
        pivot_in_0_49 <= pivot_out_0_48;
        start_in_0_49 <= start_out_0_48;
     end
  
     processor_AB AB_0_49 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_49),
       .start_in   (start_in_0_49),
       .op_in      (op_in_0_49),
       .pivot_in   (pivot_in_0_49),
       .start_out  (start_out_0_49),
       .data_out   (data_out_0_49),
       .op_out     (op_out_0_49),
       .pivot_out  (pivot_out_0_49),
       .r          (r_0_49)
     );

  // row 0, col 50

     reg start_in_0_50;
     wire start_out_0_50;

     reg [1:0] op_in_0_50;
     wire [1:0] op_out_0_50;

     wire r_0_50;

     wire data_in_0_50;
     wire data_out_0_50;

     reg pivot_in_0_50;
     wire pivot_out_0_50;

     assign data_in_0_50 = data_in[DAT_W-51];

     always @(posedge clk) begin
        op_in_0_50 <= op_out_0_49;
        pivot_in_0_50 <= pivot_out_0_49;
        start_in_0_50 <= start_out_0_49;
     end
  
     processor_AB AB_0_50 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_50),
       .start_in   (start_in_0_50),
       .op_in      (op_in_0_50),
       .pivot_in   (pivot_in_0_50),
       .start_out  (start_out_0_50),
       .data_out   (data_out_0_50),
       .op_out     (op_out_0_50),
       .pivot_out  (pivot_out_0_50),
       .r          (r_0_50)
     );

  // row 0, col 51

     reg start_in_0_51;
     wire start_out_0_51;

     reg [1:0] op_in_0_51;
     wire [1:0] op_out_0_51;

     wire r_0_51;

     wire data_in_0_51;
     wire data_out_0_51;

     reg pivot_in_0_51;
     wire pivot_out_0_51;

     assign data_in_0_51 = data_in[DAT_W-52];

     always @(posedge clk) begin
        op_in_0_51 <= op_out_0_50;
        pivot_in_0_51 <= pivot_out_0_50;
        start_in_0_51 <= start_out_0_50;
     end
  
     processor_AB AB_0_51 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_51),
       .start_in   (start_in_0_51),
       .op_in      (op_in_0_51),
       .pivot_in   (pivot_in_0_51),
       .start_out  (start_out_0_51),
       .data_out   (data_out_0_51),
       .op_out     (op_out_0_51),
       .pivot_out  (pivot_out_0_51),
       .r          (r_0_51)
     );

  // row 0, col 52

     reg start_in_0_52;
     wire start_out_0_52;

     reg [1:0] op_in_0_52;
     wire [1:0] op_out_0_52;

     wire r_0_52;

     wire data_in_0_52;
     wire data_out_0_52;

     reg pivot_in_0_52;
     wire pivot_out_0_52;

     assign data_in_0_52 = data_in[DAT_W-53];

     always @(posedge clk) begin
        op_in_0_52 <= op_out_0_51;
        pivot_in_0_52 <= pivot_out_0_51;
        start_in_0_52 <= start_out_0_51;
     end
  
     processor_AB AB_0_52 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_52),
       .start_in   (start_in_0_52),
       .op_in      (op_in_0_52),
       .pivot_in   (pivot_in_0_52),
       .start_out  (start_out_0_52),
       .data_out   (data_out_0_52),
       .op_out     (op_out_0_52),
       .pivot_out  (pivot_out_0_52),
       .r          (r_0_52)
     );

  // row 0, col 53

     reg start_in_0_53;
     wire start_out_0_53;

     reg [1:0] op_in_0_53;
     wire [1:0] op_out_0_53;

     wire r_0_53;

     wire data_in_0_53;
     wire data_out_0_53;

     reg pivot_in_0_53;
     wire pivot_out_0_53;

     assign data_in_0_53 = data_in[DAT_W-54];

     always @(posedge clk) begin
        op_in_0_53 <= op_out_0_52;
        pivot_in_0_53 <= pivot_out_0_52;
        start_in_0_53 <= start_out_0_52;
     end
  
     processor_AB AB_0_53 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_53),
       .start_in   (start_in_0_53),
       .op_in      (op_in_0_53),
       .pivot_in   (pivot_in_0_53),
       .start_out  (start_out_0_53),
       .data_out   (data_out_0_53),
       .op_out     (op_out_0_53),
       .pivot_out  (pivot_out_0_53),
       .r          (r_0_53)
     );

  // row 0, col 54

     reg start_in_0_54;
     wire start_out_0_54;

     reg [1:0] op_in_0_54;
     wire [1:0] op_out_0_54;

     wire r_0_54;

     wire data_in_0_54;
     wire data_out_0_54;

     reg pivot_in_0_54;
     wire pivot_out_0_54;

     assign data_in_0_54 = data_in[DAT_W-55];

     always @(posedge clk) begin
        op_in_0_54 <= op_out_0_53;
        pivot_in_0_54 <= pivot_out_0_53;
        start_in_0_54 <= start_out_0_53;
     end
  
     processor_AB AB_0_54 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_54),
       .start_in   (start_in_0_54),
       .op_in      (op_in_0_54),
       .pivot_in   (pivot_in_0_54),
       .start_out  (start_out_0_54),
       .data_out   (data_out_0_54),
       .op_out     (op_out_0_54),
       .pivot_out  (pivot_out_0_54),
       .r          (r_0_54)
     );

  // row 0, col 55

     reg start_in_0_55;
     wire start_out_0_55;

     reg [1:0] op_in_0_55;
     wire [1:0] op_out_0_55;

     wire r_0_55;

     wire data_in_0_55;
     wire data_out_0_55;

     reg pivot_in_0_55;
     wire pivot_out_0_55;

     assign data_in_0_55 = data_in[DAT_W-56];

     always @(posedge clk) begin
        op_in_0_55 <= op_out_0_54;
        pivot_in_0_55 <= pivot_out_0_54;
        start_in_0_55 <= start_out_0_54;
     end
  
     processor_AB AB_0_55 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_55),
       .start_in   (start_in_0_55),
       .op_in      (op_in_0_55),
       .pivot_in   (pivot_in_0_55),
       .start_out  (start_out_0_55),
       .data_out   (data_out_0_55),
       .op_out     (op_out_0_55),
       .pivot_out  (pivot_out_0_55),
       .r          (r_0_55)
     );

  // row 0, col 56

     reg start_in_0_56;
     wire start_out_0_56;

     reg [1:0] op_in_0_56;
     wire [1:0] op_out_0_56;

     wire r_0_56;

     wire data_in_0_56;
     wire data_out_0_56;

     reg pivot_in_0_56;
     wire pivot_out_0_56;

     assign data_in_0_56 = data_in[DAT_W-57];

     always @(posedge clk) begin
        op_in_0_56 <= op_out_0_55;
        pivot_in_0_56 <= pivot_out_0_55;
        start_in_0_56 <= start_out_0_55;
     end
  
     processor_AB AB_0_56 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_56),
       .start_in   (start_in_0_56),
       .op_in      (op_in_0_56),
       .pivot_in   (pivot_in_0_56),
       .start_out  (start_out_0_56),
       .data_out   (data_out_0_56),
       .op_out     (op_out_0_56),
       .pivot_out  (pivot_out_0_56),
       .r          (r_0_56)
     );

  // row 0, col 57

     reg start_in_0_57;
     wire start_out_0_57;

     reg [1:0] op_in_0_57;
     wire [1:0] op_out_0_57;

     wire r_0_57;

     wire data_in_0_57;
     wire data_out_0_57;

     reg pivot_in_0_57;
     wire pivot_out_0_57;

     assign data_in_0_57 = data_in[DAT_W-58];

     always @(posedge clk) begin
        op_in_0_57 <= op_out_0_56;
        pivot_in_0_57 <= pivot_out_0_56;
        start_in_0_57 <= start_out_0_56;
     end
  
     processor_AB AB_0_57 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_57),
       .start_in   (start_in_0_57),
       .op_in      (op_in_0_57),
       .pivot_in   (pivot_in_0_57),
       .start_out  (start_out_0_57),
       .data_out   (data_out_0_57),
       .op_out     (op_out_0_57),
       .pivot_out  (pivot_out_0_57),
       .r          (r_0_57)
     );

  // row 0, col 58

     reg start_in_0_58;
     wire start_out_0_58;

     reg [1:0] op_in_0_58;
     wire [1:0] op_out_0_58;

     wire r_0_58;

     wire data_in_0_58;
     wire data_out_0_58;

     reg pivot_in_0_58;
     wire pivot_out_0_58;

     assign data_in_0_58 = data_in[DAT_W-59];

     always @(posedge clk) begin
        op_in_0_58 <= op_out_0_57;
        pivot_in_0_58 <= pivot_out_0_57;
        start_in_0_58 <= start_out_0_57;
     end
  
     processor_AB AB_0_58 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_58),
       .start_in   (start_in_0_58),
       .op_in      (op_in_0_58),
       .pivot_in   (pivot_in_0_58),
       .start_out  (start_out_0_58),
       .data_out   (data_out_0_58),
       .op_out     (op_out_0_58),
       .pivot_out  (pivot_out_0_58),
       .r          (r_0_58)
     );

  // row 0, col 59

     reg start_in_0_59;
     wire start_out_0_59;

     reg [1:0] op_in_0_59;
     wire [1:0] op_out_0_59;

     wire r_0_59;

     wire data_in_0_59;
     wire data_out_0_59;

     reg pivot_in_0_59;
     wire pivot_out_0_59;

     assign data_in_0_59 = data_in[DAT_W-60];

     always @(posedge clk) begin
        op_in_0_59 <= op_out_0_58;
        pivot_in_0_59 <= pivot_out_0_58;
        start_in_0_59 <= start_out_0_58;
     end
  
     processor_AB AB_0_59 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_59),
       .start_in   (start_in_0_59),
       .op_in      (op_in_0_59),
       .pivot_in   (pivot_in_0_59),
       .start_out  (start_out_0_59),
       .data_out   (data_out_0_59),
       .op_out     (op_out_0_59),
       .pivot_out  (pivot_out_0_59),
       .r          (r_0_59)
     );

  // row 0, col 60

     reg start_in_0_60;
     wire start_out_0_60;

     reg [1:0] op_in_0_60;
     wire [1:0] op_out_0_60;

     wire r_0_60;

     wire data_in_0_60;
     wire data_out_0_60;

     reg pivot_in_0_60;
     wire pivot_out_0_60;

     assign data_in_0_60 = data_in[DAT_W-61];

     always @(posedge clk) begin
        op_in_0_60 <= op_out_0_59;
        pivot_in_0_60 <= pivot_out_0_59;
        start_in_0_60 <= start_out_0_59;
     end
  
     processor_AB AB_0_60 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_60),
       .start_in   (start_in_0_60),
       .op_in      (op_in_0_60),
       .pivot_in   (pivot_in_0_60),
       .start_out  (start_out_0_60),
       .data_out   (data_out_0_60),
       .op_out     (op_out_0_60),
       .pivot_out  (pivot_out_0_60),
       .r          (r_0_60)
     );

  // row 0, col 61

     reg start_in_0_61;
     wire start_out_0_61;

     reg [1:0] op_in_0_61;
     wire [1:0] op_out_0_61;

     wire r_0_61;

     wire data_in_0_61;
     wire data_out_0_61;

     reg pivot_in_0_61;
     wire pivot_out_0_61;

     assign data_in_0_61 = data_in[DAT_W-62];

     always @(posedge clk) begin
        op_in_0_61 <= op_out_0_60;
        pivot_in_0_61 <= pivot_out_0_60;
        start_in_0_61 <= start_out_0_60;
     end
  
     processor_AB AB_0_61 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_61),
       .start_in   (start_in_0_61),
       .op_in      (op_in_0_61),
       .pivot_in   (pivot_in_0_61),
       .start_out  (start_out_0_61),
       .data_out   (data_out_0_61),
       .op_out     (op_out_0_61),
       .pivot_out  (pivot_out_0_61),
       .r          (r_0_61)
     );

  // row 0, col 62

     reg start_in_0_62;
     wire start_out_0_62;

     reg [1:0] op_in_0_62;
     wire [1:0] op_out_0_62;

     wire r_0_62;

     wire data_in_0_62;
     wire data_out_0_62;

     reg pivot_in_0_62;
     wire pivot_out_0_62;

     assign data_in_0_62 = data_in[DAT_W-63];

     always @(posedge clk) begin
        op_in_0_62 <= op_out_0_61;
        pivot_in_0_62 <= pivot_out_0_61;
        start_in_0_62 <= start_out_0_61;
     end
  
     processor_AB AB_0_62 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_62),
       .start_in   (start_in_0_62),
       .op_in      (op_in_0_62),
       .pivot_in   (pivot_in_0_62),
       .start_out  (start_out_0_62),
       .data_out   (data_out_0_62),
       .op_out     (op_out_0_62),
       .pivot_out  (pivot_out_0_62),
       .r          (r_0_62)
     );

  // row 0, col 63

     reg start_in_0_63;
     wire start_out_0_63;

     reg [1:0] op_in_0_63;
     wire [1:0] op_out_0_63;

     wire r_0_63;

     wire data_in_0_63;
     wire data_out_0_63;

     reg pivot_in_0_63;
     wire pivot_out_0_63;

     assign data_in_0_63 = data_in[DAT_W-64];

     always @(posedge clk) begin
        op_in_0_63 <= op_out_0_62;
        pivot_in_0_63 <= pivot_out_0_62;
        start_in_0_63 <= start_out_0_62;
     end
  
     processor_AB AB_0_63 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_63),
       .start_in   (start_in_0_63),
       .op_in      (op_in_0_63),
       .pivot_in   (pivot_in_0_63),
       .start_out  (start_out_0_63),
       .data_out   (data_out_0_63),
       .op_out     (op_out_0_63),
       .pivot_out  (pivot_out_0_63),
       .r          (r_0_63)
     );

  // row 0, col 64

     reg start_in_0_64;
     wire start_out_0_64;

     reg [1:0] op_in_0_64;
     wire [1:0] op_out_0_64;

     wire r_0_64;

     wire data_in_0_64;
     wire data_out_0_64;

     reg pivot_in_0_64;
     wire pivot_out_0_64;

     assign data_in_0_64 = data_in[DAT_W-65];

     always @(posedge clk) begin
        op_in_0_64 <= op_out_0_63;
        pivot_in_0_64 <= pivot_out_0_63;
        start_in_0_64 <= start_out_0_63;
     end
  
     processor_AB AB_0_64 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_64),
       .start_in   (start_in_0_64),
       .op_in      (op_in_0_64),
       .pivot_in   (pivot_in_0_64),
       .start_out  (start_out_0_64),
       .data_out   (data_out_0_64),
       .op_out     (op_out_0_64),
       .pivot_out  (pivot_out_0_64),
       .r          (r_0_64)
     );

  // row 0, col 65

     reg start_in_0_65;
     wire start_out_0_65;

     reg [1:0] op_in_0_65;
     wire [1:0] op_out_0_65;

     wire r_0_65;

     wire data_in_0_65;
     wire data_out_0_65;

     reg pivot_in_0_65;
     wire pivot_out_0_65;

     assign data_in_0_65 = data_in[DAT_W-66];

     always @(posedge clk) begin
        op_in_0_65 <= op_out_0_64;
        pivot_in_0_65 <= pivot_out_0_64;
        start_in_0_65 <= start_out_0_64;
     end
  
     processor_AB AB_0_65 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_65),
       .start_in   (start_in_0_65),
       .op_in      (op_in_0_65),
       .pivot_in   (pivot_in_0_65),
       .start_out  (start_out_0_65),
       .data_out   (data_out_0_65),
       .op_out     (op_out_0_65),
       .pivot_out  (pivot_out_0_65),
       .r          (r_0_65)
     );

  // row 0, col 66

     reg start_in_0_66;
     wire start_out_0_66;

     reg [1:0] op_in_0_66;
     wire [1:0] op_out_0_66;

     wire r_0_66;

     wire data_in_0_66;
     wire data_out_0_66;

     reg pivot_in_0_66;
     wire pivot_out_0_66;

     assign data_in_0_66 = data_in[DAT_W-67];

     always @(posedge clk) begin
        op_in_0_66 <= op_out_0_65;
        pivot_in_0_66 <= pivot_out_0_65;
        start_in_0_66 <= start_out_0_65;
     end
  
     processor_AB AB_0_66 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_66),
       .start_in   (start_in_0_66),
       .op_in      (op_in_0_66),
       .pivot_in   (pivot_in_0_66),
       .start_out  (start_out_0_66),
       .data_out   (data_out_0_66),
       .op_out     (op_out_0_66),
       .pivot_out  (pivot_out_0_66),
       .r          (r_0_66)
     );

  // row 0, col 67

     reg start_in_0_67;
     wire start_out_0_67;

     reg [1:0] op_in_0_67;
     wire [1:0] op_out_0_67;

     wire r_0_67;

     wire data_in_0_67;
     wire data_out_0_67;

     reg pivot_in_0_67;
     wire pivot_out_0_67;

     assign data_in_0_67 = data_in[DAT_W-68];

     always @(posedge clk) begin
        op_in_0_67 <= op_out_0_66;
        pivot_in_0_67 <= pivot_out_0_66;
        start_in_0_67 <= start_out_0_66;
     end
  
     processor_AB AB_0_67 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_67),
       .start_in   (start_in_0_67),
       .op_in      (op_in_0_67),
       .pivot_in   (pivot_in_0_67),
       .start_out  (start_out_0_67),
       .data_out   (data_out_0_67),
       .op_out     (op_out_0_67),
       .pivot_out  (pivot_out_0_67),
       .r          (r_0_67)
     );

  // row 0, col 68

     reg start_in_0_68;
     wire start_out_0_68;

     reg [1:0] op_in_0_68;
     wire [1:0] op_out_0_68;

     wire r_0_68;

     wire data_in_0_68;
     wire data_out_0_68;

     reg pivot_in_0_68;
     wire pivot_out_0_68;

     assign data_in_0_68 = data_in[DAT_W-69];

     always @(posedge clk) begin
        op_in_0_68 <= op_out_0_67;
        pivot_in_0_68 <= pivot_out_0_67;
        start_in_0_68 <= start_out_0_67;
     end
  
     processor_AB AB_0_68 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_68),
       .start_in   (start_in_0_68),
       .op_in      (op_in_0_68),
       .pivot_in   (pivot_in_0_68),
       .start_out  (start_out_0_68),
       .data_out   (data_out_0_68),
       .op_out     (op_out_0_68),
       .pivot_out  (pivot_out_0_68),
       .r          (r_0_68)
     );

  // row 0, col 69

     reg start_in_0_69;
     wire start_out_0_69;

     reg [1:0] op_in_0_69;
     wire [1:0] op_out_0_69;

     wire r_0_69;

     wire data_in_0_69;
     wire data_out_0_69;

     reg pivot_in_0_69;
     wire pivot_out_0_69;

     assign data_in_0_69 = data_in[DAT_W-70];

     always @(posedge clk) begin
        op_in_0_69 <= op_out_0_68;
        pivot_in_0_69 <= pivot_out_0_68;
        start_in_0_69 <= start_out_0_68;
     end
  
     processor_AB AB_0_69 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_69),
       .start_in   (start_in_0_69),
       .op_in      (op_in_0_69),
       .pivot_in   (pivot_in_0_69),
       .start_out  (start_out_0_69),
       .data_out   (data_out_0_69),
       .op_out     (op_out_0_69),
       .pivot_out  (pivot_out_0_69),
       .r          (r_0_69)
     );

  // row 0, col 70

     reg start_in_0_70;
     wire start_out_0_70;

     reg [1:0] op_in_0_70;
     wire [1:0] op_out_0_70;

     wire r_0_70;

     wire data_in_0_70;
     wire data_out_0_70;

     reg pivot_in_0_70;
     wire pivot_out_0_70;

     assign data_in_0_70 = data_in[DAT_W-71];

     always @(posedge clk) begin
        op_in_0_70 <= op_out_0_69;
        pivot_in_0_70 <= pivot_out_0_69;
        start_in_0_70 <= start_out_0_69;
     end
  
     processor_AB AB_0_70 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_70),
       .start_in   (start_in_0_70),
       .op_in      (op_in_0_70),
       .pivot_in   (pivot_in_0_70),
       .start_out  (start_out_0_70),
       .data_out   (data_out_0_70),
       .op_out     (op_out_0_70),
       .pivot_out  (pivot_out_0_70),
       .r          (r_0_70)
     );

  // row 0, col 71

     reg start_in_0_71;
     wire start_out_0_71;

     reg [1:0] op_in_0_71;
     wire [1:0] op_out_0_71;

     wire r_0_71;

     wire data_in_0_71;
     wire data_out_0_71;

     reg pivot_in_0_71;
     wire pivot_out_0_71;

     assign data_in_0_71 = data_in[DAT_W-72];

     always @(posedge clk) begin
        op_in_0_71 <= op_out_0_70;
        pivot_in_0_71 <= pivot_out_0_70;
        start_in_0_71 <= start_out_0_70;
     end
  
     processor_AB AB_0_71 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_71),
       .start_in   (start_in_0_71),
       .op_in      (op_in_0_71),
       .pivot_in   (pivot_in_0_71),
       .start_out  (start_out_0_71),
       .data_out   (data_out_0_71),
       .op_out     (op_out_0_71),
       .pivot_out  (pivot_out_0_71),
       .r          (r_0_71)
     );

  // row 0, col 72

     reg start_in_0_72;
     wire start_out_0_72;

     reg [1:0] op_in_0_72;
     wire [1:0] op_out_0_72;

     wire r_0_72;

     wire data_in_0_72;
     wire data_out_0_72;

     reg pivot_in_0_72;
     wire pivot_out_0_72;

     assign data_in_0_72 = data_in[DAT_W-73];

     always @(posedge clk) begin
        op_in_0_72 <= op_out_0_71;
        pivot_in_0_72 <= pivot_out_0_71;
        start_in_0_72 <= start_out_0_71;
     end
  
     processor_AB AB_0_72 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_72),
       .start_in   (start_in_0_72),
       .op_in      (op_in_0_72),
       .pivot_in   (pivot_in_0_72),
       .start_out  (start_out_0_72),
       .data_out   (data_out_0_72),
       .op_out     (op_out_0_72),
       .pivot_out  (pivot_out_0_72),
       .r          (r_0_72)
     );

  // row 0, col 73

     reg start_in_0_73;
     wire start_out_0_73;

     reg [1:0] op_in_0_73;
     wire [1:0] op_out_0_73;

     wire r_0_73;

     wire data_in_0_73;
     wire data_out_0_73;

     reg pivot_in_0_73;
     wire pivot_out_0_73;

     assign data_in_0_73 = data_in[DAT_W-74];

     always @(posedge clk) begin
        op_in_0_73 <= op_out_0_72;
        pivot_in_0_73 <= pivot_out_0_72;
        start_in_0_73 <= start_out_0_72;
     end
  
     processor_AB AB_0_73 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_73),
       .start_in   (start_in_0_73),
       .op_in      (op_in_0_73),
       .pivot_in   (pivot_in_0_73),
       .start_out  (start_out_0_73),
       .data_out   (data_out_0_73),
       .op_out     (op_out_0_73),
       .pivot_out  (pivot_out_0_73),
       .r          (r_0_73)
     );

  // row 0, col 74

     reg start_in_0_74;
     wire start_out_0_74;

     reg [1:0] op_in_0_74;
     wire [1:0] op_out_0_74;

     wire r_0_74;

     wire data_in_0_74;
     wire data_out_0_74;

     reg pivot_in_0_74;
     wire pivot_out_0_74;

     assign data_in_0_74 = data_in[DAT_W-75];

     always @(posedge clk) begin
        op_in_0_74 <= op_out_0_73;
        pivot_in_0_74 <= pivot_out_0_73;
        start_in_0_74 <= start_out_0_73;
     end
  
     processor_AB AB_0_74 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_74),
       .start_in   (start_in_0_74),
       .op_in      (op_in_0_74),
       .pivot_in   (pivot_in_0_74),
       .start_out  (start_out_0_74),
       .data_out   (data_out_0_74),
       .op_out     (op_out_0_74),
       .pivot_out  (pivot_out_0_74),
       .r          (r_0_74)
     );

  // row 0, col 75

     reg start_in_0_75;
     wire start_out_0_75;

     reg [1:0] op_in_0_75;
     wire [1:0] op_out_0_75;

     wire r_0_75;

     wire data_in_0_75;
     wire data_out_0_75;

     reg pivot_in_0_75;
     wire pivot_out_0_75;

     assign data_in_0_75 = data_in[DAT_W-76];

     always @(posedge clk) begin
        op_in_0_75 <= op_out_0_74;
        pivot_in_0_75 <= pivot_out_0_74;
        start_in_0_75 <= start_out_0_74;
     end
  
     processor_AB AB_0_75 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_75),
       .start_in   (start_in_0_75),
       .op_in      (op_in_0_75),
       .pivot_in   (pivot_in_0_75),
       .start_out  (start_out_0_75),
       .data_out   (data_out_0_75),
       .op_out     (op_out_0_75),
       .pivot_out  (pivot_out_0_75),
       .r          (r_0_75)
     );

  // row 0, col 76

     reg start_in_0_76;
     wire start_out_0_76;

     reg [1:0] op_in_0_76;
     wire [1:0] op_out_0_76;

     wire r_0_76;

     wire data_in_0_76;
     wire data_out_0_76;

     reg pivot_in_0_76;
     wire pivot_out_0_76;

     assign data_in_0_76 = data_in[DAT_W-77];

     always @(posedge clk) begin
        op_in_0_76 <= op_out_0_75;
        pivot_in_0_76 <= pivot_out_0_75;
        start_in_0_76 <= start_out_0_75;
     end
  
     processor_AB AB_0_76 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_76),
       .start_in   (start_in_0_76),
       .op_in      (op_in_0_76),
       .pivot_in   (pivot_in_0_76),
       .start_out  (start_out_0_76),
       .data_out   (data_out_0_76),
       .op_out     (op_out_0_76),
       .pivot_out  (pivot_out_0_76),
       .r          (r_0_76)
     );

  // row 0, col 77

     reg start_in_0_77;
     wire start_out_0_77;

     reg [1:0] op_in_0_77;
     wire [1:0] op_out_0_77;

     wire r_0_77;

     wire data_in_0_77;
     wire data_out_0_77;

     reg pivot_in_0_77;
     wire pivot_out_0_77;

     assign data_in_0_77 = data_in[DAT_W-78];

     always @(posedge clk) begin
        op_in_0_77 <= op_out_0_76;
        pivot_in_0_77 <= pivot_out_0_76;
        start_in_0_77 <= start_out_0_76;
     end
  
     processor_AB AB_0_77 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_77),
       .start_in   (start_in_0_77),
       .op_in      (op_in_0_77),
       .pivot_in   (pivot_in_0_77),
       .start_out  (start_out_0_77),
       .data_out   (data_out_0_77),
       .op_out     (op_out_0_77),
       .pivot_out  (pivot_out_0_77),
       .r          (r_0_77)
     );

  // row 0, col 78

     reg start_in_0_78;
     wire start_out_0_78;

     reg [1:0] op_in_0_78;
     wire [1:0] op_out_0_78;

     wire r_0_78;

     wire data_in_0_78;
     wire data_out_0_78;

     reg pivot_in_0_78;
     wire pivot_out_0_78;

     assign data_in_0_78 = data_in[DAT_W-79];

     always @(posedge clk) begin
        op_in_0_78 <= op_out_0_77;
        pivot_in_0_78 <= pivot_out_0_77;
        start_in_0_78 <= start_out_0_77;
     end
  
     processor_AB AB_0_78 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_78),
       .start_in   (start_in_0_78),
       .op_in      (op_in_0_78),
       .pivot_in   (pivot_in_0_78),
       .start_out  (start_out_0_78),
       .data_out   (data_out_0_78),
       .op_out     (op_out_0_78),
       .pivot_out  (pivot_out_0_78),
       .r          (r_0_78)
     );

  // row 0, col 79

     reg start_in_0_79;
     wire start_out_0_79;

     reg [1:0] op_in_0_79;
     wire [1:0] op_out_0_79;

     wire r_0_79;

     wire data_in_0_79;
     wire data_out_0_79;

     reg pivot_in_0_79;
     wire pivot_out_0_79;

     assign data_in_0_79 = data_in[DAT_W-80];

     always @(posedge clk) begin
        op_in_0_79 <= op_out_0_78;
        pivot_in_0_79 <= pivot_out_0_78;
        start_in_0_79 <= start_out_0_78;
     end
  
     processor_AB AB_0_79 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_79),
       .start_in   (start_in_0_79),
       .op_in      (op_in_0_79),
       .pivot_in   (pivot_in_0_79),
       .start_out  (start_out_0_79),
       .data_out   (data_out_0_79),
       .op_out     (op_out_0_79),
       .pivot_out  (pivot_out_0_79),
       .r          (r_0_79)
     );

  // row 0, col 80

     reg start_in_0_80;
     wire start_out_0_80;

     reg [1:0] op_in_0_80;
     wire [1:0] op_out_0_80;

     wire r_0_80;

     wire data_in_0_80;
     wire data_out_0_80;

     reg pivot_in_0_80;
     wire pivot_out_0_80;

     assign data_in_0_80 = data_in[DAT_W-81];

     always @(posedge clk) begin
        op_in_0_80 <= op_out_0_79;
        pivot_in_0_80 <= pivot_out_0_79;
        start_in_0_80 <= start_out_0_79;
     end
  
     processor_AB AB_0_80 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_80),
       .start_in   (start_in_0_80),
       .op_in      (op_in_0_80),
       .pivot_in   (pivot_in_0_80),
       .start_out  (start_out_0_80),
       .data_out   (data_out_0_80),
       .op_out     (op_out_0_80),
       .pivot_out  (pivot_out_0_80),
       .r          (r_0_80)
     );

  // row 0, col 81

     reg start_in_0_81;
     wire start_out_0_81;

     reg [1:0] op_in_0_81;
     wire [1:0] op_out_0_81;

     wire r_0_81;

     wire data_in_0_81;
     wire data_out_0_81;

     reg pivot_in_0_81;
     wire pivot_out_0_81;

     assign data_in_0_81 = data_in[DAT_W-82];

     always @(posedge clk) begin
        op_in_0_81 <= op_out_0_80;
        pivot_in_0_81 <= pivot_out_0_80;
        start_in_0_81 <= start_out_0_80;
     end
  
     processor_AB AB_0_81 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_81),
       .start_in   (start_in_0_81),
       .op_in      (op_in_0_81),
       .pivot_in   (pivot_in_0_81),
       .start_out  (start_out_0_81),
       .data_out   (data_out_0_81),
       .op_out     (op_out_0_81),
       .pivot_out  (pivot_out_0_81),
       .r          (r_0_81)
     );

  // row 0, col 82

     reg start_in_0_82;
     wire start_out_0_82;

     reg [1:0] op_in_0_82;
     wire [1:0] op_out_0_82;

     wire r_0_82;

     wire data_in_0_82;
     wire data_out_0_82;

     reg pivot_in_0_82;
     wire pivot_out_0_82;

     assign data_in_0_82 = data_in[DAT_W-83];

     always @(posedge clk) begin
        op_in_0_82 <= op_out_0_81;
        pivot_in_0_82 <= pivot_out_0_81;
        start_in_0_82 <= start_out_0_81;
     end
  
     processor_AB AB_0_82 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_82),
       .start_in   (start_in_0_82),
       .op_in      (op_in_0_82),
       .pivot_in   (pivot_in_0_82),
       .start_out  (start_out_0_82),
       .data_out   (data_out_0_82),
       .op_out     (op_out_0_82),
       .pivot_out  (pivot_out_0_82),
       .r          (r_0_82)
     );

  // row 0, col 83

     reg start_in_0_83;
     wire start_out_0_83;

     reg [1:0] op_in_0_83;
     wire [1:0] op_out_0_83;

     wire r_0_83;

     wire data_in_0_83;
     wire data_out_0_83;

     reg pivot_in_0_83;
     wire pivot_out_0_83;

     assign data_in_0_83 = data_in[DAT_W-84];

     always @(posedge clk) begin
        op_in_0_83 <= op_out_0_82;
        pivot_in_0_83 <= pivot_out_0_82;
        start_in_0_83 <= start_out_0_82;
     end
  
     processor_AB AB_0_83 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_83),
       .start_in   (start_in_0_83),
       .op_in      (op_in_0_83),
       .pivot_in   (pivot_in_0_83),
       .start_out  (start_out_0_83),
       .data_out   (data_out_0_83),
       .op_out     (op_out_0_83),
       .pivot_out  (pivot_out_0_83),
       .r          (r_0_83)
     );

  // row 0, col 84

     reg start_in_0_84;
     wire start_out_0_84;

     reg [1:0] op_in_0_84;
     wire [1:0] op_out_0_84;

     wire r_0_84;

     wire data_in_0_84;
     wire data_out_0_84;

     reg pivot_in_0_84;
     wire pivot_out_0_84;

     assign data_in_0_84 = data_in[DAT_W-85];

     always @(posedge clk) begin
        op_in_0_84 <= op_out_0_83;
        pivot_in_0_84 <= pivot_out_0_83;
        start_in_0_84 <= start_out_0_83;
     end
  
     processor_AB AB_0_84 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_84),
       .start_in   (start_in_0_84),
       .op_in      (op_in_0_84),
       .pivot_in   (pivot_in_0_84),
       .start_out  (start_out_0_84),
       .data_out   (data_out_0_84),
       .op_out     (op_out_0_84),
       .pivot_out  (pivot_out_0_84),
       .r          (r_0_84)
     );

  // row 0, col 85

     reg start_in_0_85;
     wire start_out_0_85;

     reg [1:0] op_in_0_85;
     wire [1:0] op_out_0_85;

     wire r_0_85;

     wire data_in_0_85;
     wire data_out_0_85;

     reg pivot_in_0_85;
     wire pivot_out_0_85;

     assign data_in_0_85 = data_in[DAT_W-86];

     always @(posedge clk) begin
        op_in_0_85 <= op_out_0_84;
        pivot_in_0_85 <= pivot_out_0_84;
        start_in_0_85 <= start_out_0_84;
     end
  
     processor_AB AB_0_85 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_85),
       .start_in   (start_in_0_85),
       .op_in      (op_in_0_85),
       .pivot_in   (pivot_in_0_85),
       .start_out  (start_out_0_85),
       .data_out   (data_out_0_85),
       .op_out     (op_out_0_85),
       .pivot_out  (pivot_out_0_85),
       .r          (r_0_85)
     );

  // row 0, col 86

     reg start_in_0_86;
     wire start_out_0_86;

     reg [1:0] op_in_0_86;
     wire [1:0] op_out_0_86;

     wire r_0_86;

     wire data_in_0_86;
     wire data_out_0_86;

     reg pivot_in_0_86;
     wire pivot_out_0_86;

     assign data_in_0_86 = data_in[DAT_W-87];

     always @(posedge clk) begin
        op_in_0_86 <= op_out_0_85;
        pivot_in_0_86 <= pivot_out_0_85;
        start_in_0_86 <= start_out_0_85;
     end
  
     processor_AB AB_0_86 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_86),
       .start_in   (start_in_0_86),
       .op_in      (op_in_0_86),
       .pivot_in   (pivot_in_0_86),
       .start_out  (start_out_0_86),
       .data_out   (data_out_0_86),
       .op_out     (op_out_0_86),
       .pivot_out  (pivot_out_0_86),
       .r          (r_0_86)
     );

  // row 0, col 87

     reg start_in_0_87;
     wire start_out_0_87;

     reg [1:0] op_in_0_87;
     wire [1:0] op_out_0_87;

     wire r_0_87;

     wire data_in_0_87;
     wire data_out_0_87;

     reg pivot_in_0_87;
     wire pivot_out_0_87;

     assign data_in_0_87 = data_in[DAT_W-88];

     always @(posedge clk) begin
        op_in_0_87 <= op_out_0_86;
        pivot_in_0_87 <= pivot_out_0_86;
        start_in_0_87 <= start_out_0_86;
     end
  
     processor_AB AB_0_87 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_87),
       .start_in   (start_in_0_87),
       .op_in      (op_in_0_87),
       .pivot_in   (pivot_in_0_87),
       .start_out  (start_out_0_87),
       .data_out   (data_out_0_87),
       .op_out     (op_out_0_87),
       .pivot_out  (pivot_out_0_87),
       .r          (r_0_87)
     );

  // row 0, col 88

     reg start_in_0_88;
     wire start_out_0_88;

     reg [1:0] op_in_0_88;
     wire [1:0] op_out_0_88;

     wire r_0_88;

     wire data_in_0_88;
     wire data_out_0_88;

     reg pivot_in_0_88;
     wire pivot_out_0_88;

     assign data_in_0_88 = data_in[DAT_W-89];

     always @(posedge clk) begin
        op_in_0_88 <= op_out_0_87;
        pivot_in_0_88 <= pivot_out_0_87;
        start_in_0_88 <= start_out_0_87;
     end
  
     processor_AB AB_0_88 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_88),
       .start_in   (start_in_0_88),
       .op_in      (op_in_0_88),
       .pivot_in   (pivot_in_0_88),
       .start_out  (start_out_0_88),
       .data_out   (data_out_0_88),
       .op_out     (op_out_0_88),
       .pivot_out  (pivot_out_0_88),
       .r          (r_0_88)
     );

  // row 0, col 89

     reg start_in_0_89;
     wire start_out_0_89;

     reg [1:0] op_in_0_89;
     wire [1:0] op_out_0_89;

     wire r_0_89;

     wire data_in_0_89;
     wire data_out_0_89;

     reg pivot_in_0_89;
     wire pivot_out_0_89;

     assign data_in_0_89 = data_in[DAT_W-90];

     always @(posedge clk) begin
        op_in_0_89 <= op_out_0_88;
        pivot_in_0_89 <= pivot_out_0_88;
        start_in_0_89 <= start_out_0_88;
     end
  
     processor_AB AB_0_89 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_89),
       .start_in   (start_in_0_89),
       .op_in      (op_in_0_89),
       .pivot_in   (pivot_in_0_89),
       .start_out  (start_out_0_89),
       .data_out   (data_out_0_89),
       .op_out     (op_out_0_89),
       .pivot_out  (pivot_out_0_89),
       .r          (r_0_89)
     );

  // row 0, col 90

     reg start_in_0_90;
     wire start_out_0_90;

     reg [1:0] op_in_0_90;
     wire [1:0] op_out_0_90;

     wire r_0_90;

     wire data_in_0_90;
     wire data_out_0_90;

     reg pivot_in_0_90;
     wire pivot_out_0_90;

     assign data_in_0_90 = data_in[DAT_W-91];

     always @(posedge clk) begin
        op_in_0_90 <= op_out_0_89;
        pivot_in_0_90 <= pivot_out_0_89;
        start_in_0_90 <= start_out_0_89;
     end
  
     processor_AB AB_0_90 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_90),
       .start_in   (start_in_0_90),
       .op_in      (op_in_0_90),
       .pivot_in   (pivot_in_0_90),
       .start_out  (start_out_0_90),
       .data_out   (data_out_0_90),
       .op_out     (op_out_0_90),
       .pivot_out  (pivot_out_0_90),
       .r          (r_0_90)
     );

  // row 0, col 91

     reg start_in_0_91;
     wire start_out_0_91;

     reg [1:0] op_in_0_91;
     wire [1:0] op_out_0_91;

     wire r_0_91;

     wire data_in_0_91;
     wire data_out_0_91;

     reg pivot_in_0_91;
     wire pivot_out_0_91;

     assign data_in_0_91 = data_in[DAT_W-92];

     always @(posedge clk) begin
        op_in_0_91 <= op_out_0_90;
        pivot_in_0_91 <= pivot_out_0_90;
        start_in_0_91 <= start_out_0_90;
     end
  
     processor_AB AB_0_91 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_91),
       .start_in   (start_in_0_91),
       .op_in      (op_in_0_91),
       .pivot_in   (pivot_in_0_91),
       .start_out  (start_out_0_91),
       .data_out   (data_out_0_91),
       .op_out     (op_out_0_91),
       .pivot_out  (pivot_out_0_91),
       .r          (r_0_91)
     );

  // row 0, col 92

     reg start_in_0_92;
     wire start_out_0_92;

     reg [1:0] op_in_0_92;
     wire [1:0] op_out_0_92;

     wire r_0_92;

     wire data_in_0_92;
     wire data_out_0_92;

     reg pivot_in_0_92;
     wire pivot_out_0_92;

     assign data_in_0_92 = data_in[DAT_W-93];

     always @(posedge clk) begin
        op_in_0_92 <= op_out_0_91;
        pivot_in_0_92 <= pivot_out_0_91;
        start_in_0_92 <= start_out_0_91;
     end
  
     processor_AB AB_0_92 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_92),
       .start_in   (start_in_0_92),
       .op_in      (op_in_0_92),
       .pivot_in   (pivot_in_0_92),
       .start_out  (start_out_0_92),
       .data_out   (data_out_0_92),
       .op_out     (op_out_0_92),
       .pivot_out  (pivot_out_0_92),
       .r          (r_0_92)
     );

  // row 0, col 93

     reg start_in_0_93;
     wire start_out_0_93;

     reg [1:0] op_in_0_93;
     wire [1:0] op_out_0_93;

     wire r_0_93;

     wire data_in_0_93;
     wire data_out_0_93;

     reg pivot_in_0_93;
     wire pivot_out_0_93;

     assign data_in_0_93 = data_in[DAT_W-94];

     always @(posedge clk) begin
        op_in_0_93 <= op_out_0_92;
        pivot_in_0_93 <= pivot_out_0_92;
        start_in_0_93 <= start_out_0_92;
     end
  
     processor_AB AB_0_93 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_93),
       .start_in   (start_in_0_93),
       .op_in      (op_in_0_93),
       .pivot_in   (pivot_in_0_93),
       .start_out  (start_out_0_93),
       .data_out   (data_out_0_93),
       .op_out     (op_out_0_93),
       .pivot_out  (pivot_out_0_93),
       .r          (r_0_93)
     );

  // row 0, col 94

     reg start_in_0_94;
     wire start_out_0_94;

     reg [1:0] op_in_0_94;
     wire [1:0] op_out_0_94;

     wire r_0_94;

     wire data_in_0_94;
     wire data_out_0_94;

     reg pivot_in_0_94;
     wire pivot_out_0_94;

     assign data_in_0_94 = data_in[DAT_W-95];

     always @(posedge clk) begin
        op_in_0_94 <= op_out_0_93;
        pivot_in_0_94 <= pivot_out_0_93;
        start_in_0_94 <= start_out_0_93;
     end
  
     processor_AB AB_0_94 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_94),
       .start_in   (start_in_0_94),
       .op_in      (op_in_0_94),
       .pivot_in   (pivot_in_0_94),
       .start_out  (start_out_0_94),
       .data_out   (data_out_0_94),
       .op_out     (op_out_0_94),
       .pivot_out  (pivot_out_0_94),
       .r          (r_0_94)
     );

  // row 0, col 95

     reg start_in_0_95;
     wire start_out_0_95;

     reg [1:0] op_in_0_95;
     wire [1:0] op_out_0_95;

     wire r_0_95;

     wire data_in_0_95;
     wire data_out_0_95;

     reg pivot_in_0_95;
     wire pivot_out_0_95;

     assign data_in_0_95 = data_in[DAT_W-96];

     always @(posedge clk) begin
        op_in_0_95 <= op_out_0_94;
        pivot_in_0_95 <= pivot_out_0_94;
        start_in_0_95 <= start_out_0_94;
     end
  
     processor_AB AB_0_95 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_95),
       .start_in   (start_in_0_95),
       .op_in      (op_in_0_95),
       .pivot_in   (pivot_in_0_95),
       .start_out  (start_out_0_95),
       .data_out   (data_out_0_95),
       .op_out     (op_out_0_95),
       .pivot_out  (pivot_out_0_95),
       .r          (r_0_95)
     );

  // row 0, col 96

     reg start_in_0_96;
     wire start_out_0_96;

     reg [1:0] op_in_0_96;
     wire [1:0] op_out_0_96;

     wire r_0_96;

     wire data_in_0_96;
     wire data_out_0_96;

     reg pivot_in_0_96;
     wire pivot_out_0_96;

     assign data_in_0_96 = data_in[DAT_W-97];

     always @(posedge clk) begin
        op_in_0_96 <= op_out_0_95;
        pivot_in_0_96 <= pivot_out_0_95;
        start_in_0_96 <= start_out_0_95;
     end
  
     processor_AB AB_0_96 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_96),
       .start_in   (start_in_0_96),
       .op_in      (op_in_0_96),
       .pivot_in   (pivot_in_0_96),
       .start_out  (start_out_0_96),
       .data_out   (data_out_0_96),
       .op_out     (op_out_0_96),
       .pivot_out  (pivot_out_0_96),
       .r          (r_0_96)
     );

  // row 0, col 97

     reg start_in_0_97;
     wire start_out_0_97;

     reg [1:0] op_in_0_97;
     wire [1:0] op_out_0_97;

     wire r_0_97;

     wire data_in_0_97;
     wire data_out_0_97;

     reg pivot_in_0_97;
     wire pivot_out_0_97;

     assign data_in_0_97 = data_in[DAT_W-98];

     always @(posedge clk) begin
        op_in_0_97 <= op_out_0_96;
        pivot_in_0_97 <= pivot_out_0_96;
        start_in_0_97 <= start_out_0_96;
     end
  
     processor_AB AB_0_97 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_97),
       .start_in   (start_in_0_97),
       .op_in      (op_in_0_97),
       .pivot_in   (pivot_in_0_97),
       .start_out  (start_out_0_97),
       .data_out   (data_out_0_97),
       .op_out     (op_out_0_97),
       .pivot_out  (pivot_out_0_97),
       .r          (r_0_97)
     );

  // row 0, col 98

     reg start_in_0_98;
     wire start_out_0_98;

     reg [1:0] op_in_0_98;
     wire [1:0] op_out_0_98;

     wire r_0_98;

     wire data_in_0_98;
     wire data_out_0_98;

     reg pivot_in_0_98;
     wire pivot_out_0_98;

     assign data_in_0_98 = data_in[DAT_W-99];

     always @(posedge clk) begin
        op_in_0_98 <= op_out_0_97;
        pivot_in_0_98 <= pivot_out_0_97;
        start_in_0_98 <= start_out_0_97;
     end
  
     processor_AB AB_0_98 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_98),
       .start_in   (start_in_0_98),
       .op_in      (op_in_0_98),
       .pivot_in   (pivot_in_0_98),
       .start_out  (start_out_0_98),
       .data_out   (data_out_0_98),
       .op_out     (op_out_0_98),
       .pivot_out  (pivot_out_0_98),
       .r          (r_0_98)
     );

  // row 0, col 99

     reg start_in_0_99;
     wire start_out_0_99;

     reg [1:0] op_in_0_99;
     wire [1:0] op_out_0_99;

     wire r_0_99;

     wire data_in_0_99;
     wire data_out_0_99;

     reg pivot_in_0_99;
     wire pivot_out_0_99;

     assign data_in_0_99 = data_in[DAT_W-100];

     always @(posedge clk) begin
        op_in_0_99 <= op_out_0_98;
        pivot_in_0_99 <= pivot_out_0_98;
        start_in_0_99 <= start_out_0_98;
     end
  
     processor_AB AB_0_99 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_99),
       .start_in   (start_in_0_99),
       .op_in      (op_in_0_99),
       .pivot_in   (pivot_in_0_99),
       .start_out  (start_out_0_99),
       .data_out   (data_out_0_99),
       .op_out     (op_out_0_99),
       .pivot_out  (pivot_out_0_99),
       .r          (r_0_99)
     );

  // row 0, col 100

     reg start_in_0_100;
     wire start_out_0_100;

     reg [1:0] op_in_0_100;
     wire [1:0] op_out_0_100;

     wire r_0_100;

     wire data_in_0_100;
     wire data_out_0_100;

     reg pivot_in_0_100;
     wire pivot_out_0_100;

     assign data_in_0_100 = data_in[DAT_W-101];

     always @(posedge clk) begin
        op_in_0_100 <= op_out_0_99;
        pivot_in_0_100 <= pivot_out_0_99;
        start_in_0_100 <= start_out_0_99;
     end
  
     processor_AB AB_0_100 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_100),
       .start_in   (start_in_0_100),
       .op_in      (op_in_0_100),
       .pivot_in   (pivot_in_0_100),
       .start_out  (start_out_0_100),
       .data_out   (data_out_0_100),
       .op_out     (op_out_0_100),
       .pivot_out  (pivot_out_0_100),
       .r          (r_0_100)
     );

  /////////////////////////////////////
  // row 1
  // row 1, col 0

     wire start_in_1_0;
     wire start_out_1_0;

     wire [1:0] op_in_1_0;
     wire [1:0] op_out_1_0;

     wire r_1_0;

     reg data_in_1_0;
     wire data_out_1_0;

     wire pivot_in_1_0;
     wire pivout_out_1_0;

     assign op_in_1_0 = mode & start ? 2'b01 : 2'b00;
     assign pivot_in_1_0 = 0;

     assign start_in_1_0 = start_row[1]; 

     always @(posedge clk) begin
         data_in_1_0 <= data_out_0_0;
     end

     processor_AB AB_1_0 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_0),
       .start_in   (start_in_1_0),
       .op_in      (op_in_1_0),
       .pivot_in   (pivot_in_1_0),
       .start_out  (start_out_1_0),
       .data_out   (data_out_1_0),
       .op_out     (op_out_1_0),
       .pivot_out  (pivot_out_1_0),
       .r          (r_1_0)
     );

  // row 1, col 1

     reg start_in_1_1;
     wire start_out_1_1;

     reg [1:0] op_in_1_1;
     wire [1:0] op_out_1_1;

     wire r_1_1;

     reg data_in_1_1;
     wire data_out_1_1;

     reg pivot_in_1_1;
     wire pivot_out_1_1;

     always @(posedge clk) begin
         op_in_1_1 <= op_out_1_0;
         pivot_in_1_1 <= pivot_out_1_0;
         start_in_1_1 <= start_out_1_0;
     end

     always @(posedge clk) begin
         data_in_1_1 <= data_out_0_1;
     end
  
     processor_AB AB_1_1 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_1),
       .start_in   (start_in_1_1),
       .op_in      (op_in_1_1),
       .pivot_in   (pivot_in_1_1),
       .start_out  (start_out_1_1),
       .data_out   (data_out_1_1),
       .op_out     (op_out_1_1),
       .pivot_out  (pivot_out_1_1),
       .r          (r_1_1)
     );

  // row 1, col 2

     reg start_in_1_2;
     wire start_out_1_2;

     reg [1:0] op_in_1_2;
     wire [1:0] op_out_1_2;

     wire r_1_2;

     reg data_in_1_2;
     wire data_out_1_2;

     reg pivot_in_1_2;
     wire pivot_out_1_2;

     always @(posedge clk) begin
         op_in_1_2 <= op_out_1_1;
         pivot_in_1_2 <= pivot_out_1_1;
         start_in_1_2 <= start_out_1_1;
     end

     always @(posedge clk) begin
         data_in_1_2 <= data_out_0_2;
     end
  
     processor_AB AB_1_2 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_2),
       .start_in   (start_in_1_2),
       .op_in      (op_in_1_2),
       .pivot_in   (pivot_in_1_2),
       .start_out  (start_out_1_2),
       .data_out   (data_out_1_2),
       .op_out     (op_out_1_2),
       .pivot_out  (pivot_out_1_2),
       .r          (r_1_2)
     );

  // row 1, col 3

     reg start_in_1_3;
     wire start_out_1_3;

     reg [1:0] op_in_1_3;
     wire [1:0] op_out_1_3;

     wire r_1_3;

     reg data_in_1_3;
     wire data_out_1_3;

     reg pivot_in_1_3;
     wire pivot_out_1_3;

     always @(posedge clk) begin
         op_in_1_3 <= op_out_1_2;
         pivot_in_1_3 <= pivot_out_1_2;
         start_in_1_3 <= start_out_1_2;
     end

     always @(posedge clk) begin
         data_in_1_3 <= data_out_0_3;
     end
  
     processor_AB AB_1_3 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_3),
       .start_in   (start_in_1_3),
       .op_in      (op_in_1_3),
       .pivot_in   (pivot_in_1_3),
       .start_out  (start_out_1_3),
       .data_out   (data_out_1_3),
       .op_out     (op_out_1_3),
       .pivot_out  (pivot_out_1_3),
       .r          (r_1_3)
     );

  // row 1, col 4

     reg start_in_1_4;
     wire start_out_1_4;

     reg [1:0] op_in_1_4;
     wire [1:0] op_out_1_4;

     wire r_1_4;

     reg data_in_1_4;
     wire data_out_1_4;

     reg pivot_in_1_4;
     wire pivot_out_1_4;

     always @(posedge clk) begin
         op_in_1_4 <= op_out_1_3;
         pivot_in_1_4 <= pivot_out_1_3;
         start_in_1_4 <= start_out_1_3;
     end

     always @(posedge clk) begin
         data_in_1_4 <= data_out_0_4;
     end
  
     processor_AB AB_1_4 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_4),
       .start_in   (start_in_1_4),
       .op_in      (op_in_1_4),
       .pivot_in   (pivot_in_1_4),
       .start_out  (start_out_1_4),
       .data_out   (data_out_1_4),
       .op_out     (op_out_1_4),
       .pivot_out  (pivot_out_1_4),
       .r          (r_1_4)
     );

  // row 1, col 5

     reg start_in_1_5;
     wire start_out_1_5;

     reg [1:0] op_in_1_5;
     wire [1:0] op_out_1_5;

     wire r_1_5;

     reg data_in_1_5;
     wire data_out_1_5;

     reg pivot_in_1_5;
     wire pivot_out_1_5;

     always @(posedge clk) begin
         op_in_1_5 <= op_out_1_4;
         pivot_in_1_5 <= pivot_out_1_4;
         start_in_1_5 <= start_out_1_4;
     end

     always @(posedge clk) begin
         data_in_1_5 <= data_out_0_5;
     end
  
     processor_AB AB_1_5 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_5),
       .start_in   (start_in_1_5),
       .op_in      (op_in_1_5),
       .pivot_in   (pivot_in_1_5),
       .start_out  (start_out_1_5),
       .data_out   (data_out_1_5),
       .op_out     (op_out_1_5),
       .pivot_out  (pivot_out_1_5),
       .r          (r_1_5)
     );

  // row 1, col 6

     reg start_in_1_6;
     wire start_out_1_6;

     reg [1:0] op_in_1_6;
     wire [1:0] op_out_1_6;

     wire r_1_6;

     reg data_in_1_6;
     wire data_out_1_6;

     reg pivot_in_1_6;
     wire pivot_out_1_6;

     always @(posedge clk) begin
         op_in_1_6 <= op_out_1_5;
         pivot_in_1_6 <= pivot_out_1_5;
         start_in_1_6 <= start_out_1_5;
     end

     always @(posedge clk) begin
         data_in_1_6 <= data_out_0_6;
     end
  
     processor_AB AB_1_6 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_6),
       .start_in   (start_in_1_6),
       .op_in      (op_in_1_6),
       .pivot_in   (pivot_in_1_6),
       .start_out  (start_out_1_6),
       .data_out   (data_out_1_6),
       .op_out     (op_out_1_6),
       .pivot_out  (pivot_out_1_6),
       .r          (r_1_6)
     );

  // row 1, col 7

     reg start_in_1_7;
     wire start_out_1_7;

     reg [1:0] op_in_1_7;
     wire [1:0] op_out_1_7;

     wire r_1_7;

     reg data_in_1_7;
     wire data_out_1_7;

     reg pivot_in_1_7;
     wire pivot_out_1_7;

     always @(posedge clk) begin
         op_in_1_7 <= op_out_1_6;
         pivot_in_1_7 <= pivot_out_1_6;
         start_in_1_7 <= start_out_1_6;
     end

     always @(posedge clk) begin
         data_in_1_7 <= data_out_0_7;
     end
  
     processor_AB AB_1_7 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_7),
       .start_in   (start_in_1_7),
       .op_in      (op_in_1_7),
       .pivot_in   (pivot_in_1_7),
       .start_out  (start_out_1_7),
       .data_out   (data_out_1_7),
       .op_out     (op_out_1_7),
       .pivot_out  (pivot_out_1_7),
       .r          (r_1_7)
     );

  // row 1, col 8

     reg start_in_1_8;
     wire start_out_1_8;

     reg [1:0] op_in_1_8;
     wire [1:0] op_out_1_8;

     wire r_1_8;

     reg data_in_1_8;
     wire data_out_1_8;

     reg pivot_in_1_8;
     wire pivot_out_1_8;

     always @(posedge clk) begin
         op_in_1_8 <= op_out_1_7;
         pivot_in_1_8 <= pivot_out_1_7;
         start_in_1_8 <= start_out_1_7;
     end

     always @(posedge clk) begin
         data_in_1_8 <= data_out_0_8;
     end
  
     processor_AB AB_1_8 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_8),
       .start_in   (start_in_1_8),
       .op_in      (op_in_1_8),
       .pivot_in   (pivot_in_1_8),
       .start_out  (start_out_1_8),
       .data_out   (data_out_1_8),
       .op_out     (op_out_1_8),
       .pivot_out  (pivot_out_1_8),
       .r          (r_1_8)
     );

  // row 1, col 9

     reg start_in_1_9;
     wire start_out_1_9;

     reg [1:0] op_in_1_9;
     wire [1:0] op_out_1_9;

     wire r_1_9;

     reg data_in_1_9;
     wire data_out_1_9;

     reg pivot_in_1_9;
     wire pivot_out_1_9;

     always @(posedge clk) begin
         op_in_1_9 <= op_out_1_8;
         pivot_in_1_9 <= pivot_out_1_8;
         start_in_1_9 <= start_out_1_8;
     end

     always @(posedge clk) begin
         data_in_1_9 <= data_out_0_9;
     end
  
     processor_AB AB_1_9 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_9),
       .start_in   (start_in_1_9),
       .op_in      (op_in_1_9),
       .pivot_in   (pivot_in_1_9),
       .start_out  (start_out_1_9),
       .data_out   (data_out_1_9),
       .op_out     (op_out_1_9),
       .pivot_out  (pivot_out_1_9),
       .r          (r_1_9)
     );

  // row 1, col 10

     reg start_in_1_10;
     wire start_out_1_10;

     reg [1:0] op_in_1_10;
     wire [1:0] op_out_1_10;

     wire r_1_10;

     reg data_in_1_10;
     wire data_out_1_10;

     reg pivot_in_1_10;
     wire pivot_out_1_10;

     always @(posedge clk) begin
         op_in_1_10 <= op_out_1_9;
         pivot_in_1_10 <= pivot_out_1_9;
         start_in_1_10 <= start_out_1_9;
     end

     always @(posedge clk) begin
         data_in_1_10 <= data_out_0_10;
     end
  
     processor_AB AB_1_10 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_10),
       .start_in   (start_in_1_10),
       .op_in      (op_in_1_10),
       .pivot_in   (pivot_in_1_10),
       .start_out  (start_out_1_10),
       .data_out   (data_out_1_10),
       .op_out     (op_out_1_10),
       .pivot_out  (pivot_out_1_10),
       .r          (r_1_10)
     );

  // row 1, col 11

     reg start_in_1_11;
     wire start_out_1_11;

     reg [1:0] op_in_1_11;
     wire [1:0] op_out_1_11;

     wire r_1_11;

     reg data_in_1_11;
     wire data_out_1_11;

     reg pivot_in_1_11;
     wire pivot_out_1_11;

     always @(posedge clk) begin
         op_in_1_11 <= op_out_1_10;
         pivot_in_1_11 <= pivot_out_1_10;
         start_in_1_11 <= start_out_1_10;
     end

     always @(posedge clk) begin
         data_in_1_11 <= data_out_0_11;
     end
  
     processor_AB AB_1_11 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_11),
       .start_in   (start_in_1_11),
       .op_in      (op_in_1_11),
       .pivot_in   (pivot_in_1_11),
       .start_out  (start_out_1_11),
       .data_out   (data_out_1_11),
       .op_out     (op_out_1_11),
       .pivot_out  (pivot_out_1_11),
       .r          (r_1_11)
     );

  // row 1, col 12

     reg start_in_1_12;
     wire start_out_1_12;

     reg [1:0] op_in_1_12;
     wire [1:0] op_out_1_12;

     wire r_1_12;

     reg data_in_1_12;
     wire data_out_1_12;

     reg pivot_in_1_12;
     wire pivot_out_1_12;

     always @(posedge clk) begin
         op_in_1_12 <= op_out_1_11;
         pivot_in_1_12 <= pivot_out_1_11;
         start_in_1_12 <= start_out_1_11;
     end

     always @(posedge clk) begin
         data_in_1_12 <= data_out_0_12;
     end
  
     processor_AB AB_1_12 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_12),
       .start_in   (start_in_1_12),
       .op_in      (op_in_1_12),
       .pivot_in   (pivot_in_1_12),
       .start_out  (start_out_1_12),
       .data_out   (data_out_1_12),
       .op_out     (op_out_1_12),
       .pivot_out  (pivot_out_1_12),
       .r          (r_1_12)
     );

  // row 1, col 13

     reg start_in_1_13;
     wire start_out_1_13;

     reg [1:0] op_in_1_13;
     wire [1:0] op_out_1_13;

     wire r_1_13;

     reg data_in_1_13;
     wire data_out_1_13;

     reg pivot_in_1_13;
     wire pivot_out_1_13;

     always @(posedge clk) begin
         op_in_1_13 <= op_out_1_12;
         pivot_in_1_13 <= pivot_out_1_12;
         start_in_1_13 <= start_out_1_12;
     end

     always @(posedge clk) begin
         data_in_1_13 <= data_out_0_13;
     end
  
     processor_AB AB_1_13 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_13),
       .start_in   (start_in_1_13),
       .op_in      (op_in_1_13),
       .pivot_in   (pivot_in_1_13),
       .start_out  (start_out_1_13),
       .data_out   (data_out_1_13),
       .op_out     (op_out_1_13),
       .pivot_out  (pivot_out_1_13),
       .r          (r_1_13)
     );

  // row 1, col 14

     reg start_in_1_14;
     wire start_out_1_14;

     reg [1:0] op_in_1_14;
     wire [1:0] op_out_1_14;

     wire r_1_14;

     reg data_in_1_14;
     wire data_out_1_14;

     reg pivot_in_1_14;
     wire pivot_out_1_14;

     always @(posedge clk) begin
         op_in_1_14 <= op_out_1_13;
         pivot_in_1_14 <= pivot_out_1_13;
         start_in_1_14 <= start_out_1_13;
     end

     always @(posedge clk) begin
         data_in_1_14 <= data_out_0_14;
     end
  
     processor_AB AB_1_14 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_14),
       .start_in   (start_in_1_14),
       .op_in      (op_in_1_14),
       .pivot_in   (pivot_in_1_14),
       .start_out  (start_out_1_14),
       .data_out   (data_out_1_14),
       .op_out     (op_out_1_14),
       .pivot_out  (pivot_out_1_14),
       .r          (r_1_14)
     );

  // row 1, col 15

     reg start_in_1_15;
     wire start_out_1_15;

     reg [1:0] op_in_1_15;
     wire [1:0] op_out_1_15;

     wire r_1_15;

     reg data_in_1_15;
     wire data_out_1_15;

     reg pivot_in_1_15;
     wire pivot_out_1_15;

     always @(posedge clk) begin
         op_in_1_15 <= op_out_1_14;
         pivot_in_1_15 <= pivot_out_1_14;
         start_in_1_15 <= start_out_1_14;
     end

     always @(posedge clk) begin
         data_in_1_15 <= data_out_0_15;
     end
  
     processor_AB AB_1_15 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_15),
       .start_in   (start_in_1_15),
       .op_in      (op_in_1_15),
       .pivot_in   (pivot_in_1_15),
       .start_out  (start_out_1_15),
       .data_out   (data_out_1_15),
       .op_out     (op_out_1_15),
       .pivot_out  (pivot_out_1_15),
       .r          (r_1_15)
     );

  // row 1, col 16

     reg start_in_1_16;
     wire start_out_1_16;

     reg [1:0] op_in_1_16;
     wire [1:0] op_out_1_16;

     wire r_1_16;

     reg data_in_1_16;
     wire data_out_1_16;

     reg pivot_in_1_16;
     wire pivot_out_1_16;

     always @(posedge clk) begin
         op_in_1_16 <= op_out_1_15;
         pivot_in_1_16 <= pivot_out_1_15;
         start_in_1_16 <= start_out_1_15;
     end

     always @(posedge clk) begin
         data_in_1_16 <= data_out_0_16;
     end
  
     processor_AB AB_1_16 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_16),
       .start_in   (start_in_1_16),
       .op_in      (op_in_1_16),
       .pivot_in   (pivot_in_1_16),
       .start_out  (start_out_1_16),
       .data_out   (data_out_1_16),
       .op_out     (op_out_1_16),
       .pivot_out  (pivot_out_1_16),
       .r          (r_1_16)
     );

  // row 1, col 17

     reg start_in_1_17;
     wire start_out_1_17;

     reg [1:0] op_in_1_17;
     wire [1:0] op_out_1_17;

     wire r_1_17;

     reg data_in_1_17;
     wire data_out_1_17;

     reg pivot_in_1_17;
     wire pivot_out_1_17;

     always @(posedge clk) begin
         op_in_1_17 <= op_out_1_16;
         pivot_in_1_17 <= pivot_out_1_16;
         start_in_1_17 <= start_out_1_16;
     end

     always @(posedge clk) begin
         data_in_1_17 <= data_out_0_17;
     end
  
     processor_AB AB_1_17 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_17),
       .start_in   (start_in_1_17),
       .op_in      (op_in_1_17),
       .pivot_in   (pivot_in_1_17),
       .start_out  (start_out_1_17),
       .data_out   (data_out_1_17),
       .op_out     (op_out_1_17),
       .pivot_out  (pivot_out_1_17),
       .r          (r_1_17)
     );

  // row 1, col 18

     reg start_in_1_18;
     wire start_out_1_18;

     reg [1:0] op_in_1_18;
     wire [1:0] op_out_1_18;

     wire r_1_18;

     reg data_in_1_18;
     wire data_out_1_18;

     reg pivot_in_1_18;
     wire pivot_out_1_18;

     always @(posedge clk) begin
         op_in_1_18 <= op_out_1_17;
         pivot_in_1_18 <= pivot_out_1_17;
         start_in_1_18 <= start_out_1_17;
     end

     always @(posedge clk) begin
         data_in_1_18 <= data_out_0_18;
     end
  
     processor_AB AB_1_18 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_18),
       .start_in   (start_in_1_18),
       .op_in      (op_in_1_18),
       .pivot_in   (pivot_in_1_18),
       .start_out  (start_out_1_18),
       .data_out   (data_out_1_18),
       .op_out     (op_out_1_18),
       .pivot_out  (pivot_out_1_18),
       .r          (r_1_18)
     );

  // row 1, col 19

     reg start_in_1_19;
     wire start_out_1_19;

     reg [1:0] op_in_1_19;
     wire [1:0] op_out_1_19;

     wire r_1_19;

     reg data_in_1_19;
     wire data_out_1_19;

     reg pivot_in_1_19;
     wire pivot_out_1_19;

     always @(posedge clk) begin
         op_in_1_19 <= op_out_1_18;
         pivot_in_1_19 <= pivot_out_1_18;
         start_in_1_19 <= start_out_1_18;
     end

     always @(posedge clk) begin
         data_in_1_19 <= data_out_0_19;
     end
  
     processor_AB AB_1_19 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_19),
       .start_in   (start_in_1_19),
       .op_in      (op_in_1_19),
       .pivot_in   (pivot_in_1_19),
       .start_out  (start_out_1_19),
       .data_out   (data_out_1_19),
       .op_out     (op_out_1_19),
       .pivot_out  (pivot_out_1_19),
       .r          (r_1_19)
     );

  // row 1, col 20

     reg start_in_1_20;
     wire start_out_1_20;

     reg [1:0] op_in_1_20;
     wire [1:0] op_out_1_20;

     wire r_1_20;

     reg data_in_1_20;
     wire data_out_1_20;

     reg pivot_in_1_20;
     wire pivot_out_1_20;

     always @(posedge clk) begin
         op_in_1_20 <= op_out_1_19;
         pivot_in_1_20 <= pivot_out_1_19;
         start_in_1_20 <= start_out_1_19;
     end

     always @(posedge clk) begin
         data_in_1_20 <= data_out_0_20;
     end
  
     processor_AB AB_1_20 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_20),
       .start_in   (start_in_1_20),
       .op_in      (op_in_1_20),
       .pivot_in   (pivot_in_1_20),
       .start_out  (start_out_1_20),
       .data_out   (data_out_1_20),
       .op_out     (op_out_1_20),
       .pivot_out  (pivot_out_1_20),
       .r          (r_1_20)
     );

  // row 1, col 21

     reg start_in_1_21;
     wire start_out_1_21;

     reg [1:0] op_in_1_21;
     wire [1:0] op_out_1_21;

     wire r_1_21;

     reg data_in_1_21;
     wire data_out_1_21;

     reg pivot_in_1_21;
     wire pivot_out_1_21;

     always @(posedge clk) begin
         op_in_1_21 <= op_out_1_20;
         pivot_in_1_21 <= pivot_out_1_20;
         start_in_1_21 <= start_out_1_20;
     end

     always @(posedge clk) begin
         data_in_1_21 <= data_out_0_21;
     end
  
     processor_AB AB_1_21 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_21),
       .start_in   (start_in_1_21),
       .op_in      (op_in_1_21),
       .pivot_in   (pivot_in_1_21),
       .start_out  (start_out_1_21),
       .data_out   (data_out_1_21),
       .op_out     (op_out_1_21),
       .pivot_out  (pivot_out_1_21),
       .r          (r_1_21)
     );

  // row 1, col 22

     reg start_in_1_22;
     wire start_out_1_22;

     reg [1:0] op_in_1_22;
     wire [1:0] op_out_1_22;

     wire r_1_22;

     reg data_in_1_22;
     wire data_out_1_22;

     reg pivot_in_1_22;
     wire pivot_out_1_22;

     always @(posedge clk) begin
         op_in_1_22 <= op_out_1_21;
         pivot_in_1_22 <= pivot_out_1_21;
         start_in_1_22 <= start_out_1_21;
     end

     always @(posedge clk) begin
         data_in_1_22 <= data_out_0_22;
     end
  
     processor_AB AB_1_22 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_22),
       .start_in   (start_in_1_22),
       .op_in      (op_in_1_22),
       .pivot_in   (pivot_in_1_22),
       .start_out  (start_out_1_22),
       .data_out   (data_out_1_22),
       .op_out     (op_out_1_22),
       .pivot_out  (pivot_out_1_22),
       .r          (r_1_22)
     );

  // row 1, col 23

     reg start_in_1_23;
     wire start_out_1_23;

     reg [1:0] op_in_1_23;
     wire [1:0] op_out_1_23;

     wire r_1_23;

     reg data_in_1_23;
     wire data_out_1_23;

     reg pivot_in_1_23;
     wire pivot_out_1_23;

     always @(posedge clk) begin
         op_in_1_23 <= op_out_1_22;
         pivot_in_1_23 <= pivot_out_1_22;
         start_in_1_23 <= start_out_1_22;
     end

     always @(posedge clk) begin
         data_in_1_23 <= data_out_0_23;
     end
  
     processor_AB AB_1_23 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_23),
       .start_in   (start_in_1_23),
       .op_in      (op_in_1_23),
       .pivot_in   (pivot_in_1_23),
       .start_out  (start_out_1_23),
       .data_out   (data_out_1_23),
       .op_out     (op_out_1_23),
       .pivot_out  (pivot_out_1_23),
       .r          (r_1_23)
     );

  // row 1, col 24

     reg start_in_1_24;
     wire start_out_1_24;

     reg [1:0] op_in_1_24;
     wire [1:0] op_out_1_24;

     wire r_1_24;

     reg data_in_1_24;
     wire data_out_1_24;

     reg pivot_in_1_24;
     wire pivot_out_1_24;

     always @(posedge clk) begin
         op_in_1_24 <= op_out_1_23;
         pivot_in_1_24 <= pivot_out_1_23;
         start_in_1_24 <= start_out_1_23;
     end

     always @(posedge clk) begin
         data_in_1_24 <= data_out_0_24;
     end
  
     processor_AB AB_1_24 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_24),
       .start_in   (start_in_1_24),
       .op_in      (op_in_1_24),
       .pivot_in   (pivot_in_1_24),
       .start_out  (start_out_1_24),
       .data_out   (data_out_1_24),
       .op_out     (op_out_1_24),
       .pivot_out  (pivot_out_1_24),
       .r          (r_1_24)
     );

  // row 1, col 25

     reg start_in_1_25;
     wire start_out_1_25;

     reg [1:0] op_in_1_25;
     wire [1:0] op_out_1_25;

     wire r_1_25;

     reg data_in_1_25;
     wire data_out_1_25;

     reg pivot_in_1_25;
     wire pivot_out_1_25;

     always @(posedge clk) begin
         op_in_1_25 <= op_out_1_24;
         pivot_in_1_25 <= pivot_out_1_24;
         start_in_1_25 <= start_out_1_24;
     end

     always @(posedge clk) begin
         data_in_1_25 <= data_out_0_25;
     end
  
     processor_AB AB_1_25 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_25),
       .start_in   (start_in_1_25),
       .op_in      (op_in_1_25),
       .pivot_in   (pivot_in_1_25),
       .start_out  (start_out_1_25),
       .data_out   (data_out_1_25),
       .op_out     (op_out_1_25),
       .pivot_out  (pivot_out_1_25),
       .r          (r_1_25)
     );

  // row 1, col 26

     reg start_in_1_26;
     wire start_out_1_26;

     reg [1:0] op_in_1_26;
     wire [1:0] op_out_1_26;

     wire r_1_26;

     reg data_in_1_26;
     wire data_out_1_26;

     reg pivot_in_1_26;
     wire pivot_out_1_26;

     always @(posedge clk) begin
         op_in_1_26 <= op_out_1_25;
         pivot_in_1_26 <= pivot_out_1_25;
         start_in_1_26 <= start_out_1_25;
     end

     always @(posedge clk) begin
         data_in_1_26 <= data_out_0_26;
     end
  
     processor_AB AB_1_26 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_26),
       .start_in   (start_in_1_26),
       .op_in      (op_in_1_26),
       .pivot_in   (pivot_in_1_26),
       .start_out  (start_out_1_26),
       .data_out   (data_out_1_26),
       .op_out     (op_out_1_26),
       .pivot_out  (pivot_out_1_26),
       .r          (r_1_26)
     );

  // row 1, col 27

     reg start_in_1_27;
     wire start_out_1_27;

     reg [1:0] op_in_1_27;
     wire [1:0] op_out_1_27;

     wire r_1_27;

     reg data_in_1_27;
     wire data_out_1_27;

     reg pivot_in_1_27;
     wire pivot_out_1_27;

     always @(posedge clk) begin
         op_in_1_27 <= op_out_1_26;
         pivot_in_1_27 <= pivot_out_1_26;
         start_in_1_27 <= start_out_1_26;
     end

     always @(posedge clk) begin
         data_in_1_27 <= data_out_0_27;
     end
  
     processor_AB AB_1_27 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_27),
       .start_in   (start_in_1_27),
       .op_in      (op_in_1_27),
       .pivot_in   (pivot_in_1_27),
       .start_out  (start_out_1_27),
       .data_out   (data_out_1_27),
       .op_out     (op_out_1_27),
       .pivot_out  (pivot_out_1_27),
       .r          (r_1_27)
     );

  // row 1, col 28

     reg start_in_1_28;
     wire start_out_1_28;

     reg [1:0] op_in_1_28;
     wire [1:0] op_out_1_28;

     wire r_1_28;

     reg data_in_1_28;
     wire data_out_1_28;

     reg pivot_in_1_28;
     wire pivot_out_1_28;

     always @(posedge clk) begin
         op_in_1_28 <= op_out_1_27;
         pivot_in_1_28 <= pivot_out_1_27;
         start_in_1_28 <= start_out_1_27;
     end

     always @(posedge clk) begin
         data_in_1_28 <= data_out_0_28;
     end
  
     processor_AB AB_1_28 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_28),
       .start_in   (start_in_1_28),
       .op_in      (op_in_1_28),
       .pivot_in   (pivot_in_1_28),
       .start_out  (start_out_1_28),
       .data_out   (data_out_1_28),
       .op_out     (op_out_1_28),
       .pivot_out  (pivot_out_1_28),
       .r          (r_1_28)
     );

  // row 1, col 29

     reg start_in_1_29;
     wire start_out_1_29;

     reg [1:0] op_in_1_29;
     wire [1:0] op_out_1_29;

     wire r_1_29;

     reg data_in_1_29;
     wire data_out_1_29;

     reg pivot_in_1_29;
     wire pivot_out_1_29;

     always @(posedge clk) begin
         op_in_1_29 <= op_out_1_28;
         pivot_in_1_29 <= pivot_out_1_28;
         start_in_1_29 <= start_out_1_28;
     end

     always @(posedge clk) begin
         data_in_1_29 <= data_out_0_29;
     end
  
     processor_AB AB_1_29 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_29),
       .start_in   (start_in_1_29),
       .op_in      (op_in_1_29),
       .pivot_in   (pivot_in_1_29),
       .start_out  (start_out_1_29),
       .data_out   (data_out_1_29),
       .op_out     (op_out_1_29),
       .pivot_out  (pivot_out_1_29),
       .r          (r_1_29)
     );

  // row 1, col 30

     reg start_in_1_30;
     wire start_out_1_30;

     reg [1:0] op_in_1_30;
     wire [1:0] op_out_1_30;

     wire r_1_30;

     reg data_in_1_30;
     wire data_out_1_30;

     reg pivot_in_1_30;
     wire pivot_out_1_30;

     always @(posedge clk) begin
         op_in_1_30 <= op_out_1_29;
         pivot_in_1_30 <= pivot_out_1_29;
         start_in_1_30 <= start_out_1_29;
     end

     always @(posedge clk) begin
         data_in_1_30 <= data_out_0_30;
     end
  
     processor_AB AB_1_30 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_30),
       .start_in   (start_in_1_30),
       .op_in      (op_in_1_30),
       .pivot_in   (pivot_in_1_30),
       .start_out  (start_out_1_30),
       .data_out   (data_out_1_30),
       .op_out     (op_out_1_30),
       .pivot_out  (pivot_out_1_30),
       .r          (r_1_30)
     );

  // row 1, col 31

     reg start_in_1_31;
     wire start_out_1_31;

     reg [1:0] op_in_1_31;
     wire [1:0] op_out_1_31;

     wire r_1_31;

     reg data_in_1_31;
     wire data_out_1_31;

     reg pivot_in_1_31;
     wire pivot_out_1_31;

     always @(posedge clk) begin
         op_in_1_31 <= op_out_1_30;
         pivot_in_1_31 <= pivot_out_1_30;
         start_in_1_31 <= start_out_1_30;
     end

     always @(posedge clk) begin
         data_in_1_31 <= data_out_0_31;
     end
  
     processor_AB AB_1_31 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_31),
       .start_in   (start_in_1_31),
       .op_in      (op_in_1_31),
       .pivot_in   (pivot_in_1_31),
       .start_out  (start_out_1_31),
       .data_out   (data_out_1_31),
       .op_out     (op_out_1_31),
       .pivot_out  (pivot_out_1_31),
       .r          (r_1_31)
     );

  // row 1, col 32

     reg start_in_1_32;
     wire start_out_1_32;

     reg [1:0] op_in_1_32;
     wire [1:0] op_out_1_32;

     wire r_1_32;

     reg data_in_1_32;
     wire data_out_1_32;

     reg pivot_in_1_32;
     wire pivot_out_1_32;

     always @(posedge clk) begin
         op_in_1_32 <= op_out_1_31;
         pivot_in_1_32 <= pivot_out_1_31;
         start_in_1_32 <= start_out_1_31;
     end

     always @(posedge clk) begin
         data_in_1_32 <= data_out_0_32;
     end
  
     processor_AB AB_1_32 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_32),
       .start_in   (start_in_1_32),
       .op_in      (op_in_1_32),
       .pivot_in   (pivot_in_1_32),
       .start_out  (start_out_1_32),
       .data_out   (data_out_1_32),
       .op_out     (op_out_1_32),
       .pivot_out  (pivot_out_1_32),
       .r          (r_1_32)
     );

  // row 1, col 33

     reg start_in_1_33;
     wire start_out_1_33;

     reg [1:0] op_in_1_33;
     wire [1:0] op_out_1_33;

     wire r_1_33;

     reg data_in_1_33;
     wire data_out_1_33;

     reg pivot_in_1_33;
     wire pivot_out_1_33;

     always @(posedge clk) begin
         op_in_1_33 <= op_out_1_32;
         pivot_in_1_33 <= pivot_out_1_32;
         start_in_1_33 <= start_out_1_32;
     end

     always @(posedge clk) begin
         data_in_1_33 <= data_out_0_33;
     end
  
     processor_AB AB_1_33 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_33),
       .start_in   (start_in_1_33),
       .op_in      (op_in_1_33),
       .pivot_in   (pivot_in_1_33),
       .start_out  (start_out_1_33),
       .data_out   (data_out_1_33),
       .op_out     (op_out_1_33),
       .pivot_out  (pivot_out_1_33),
       .r          (r_1_33)
     );

  // row 1, col 34

     reg start_in_1_34;
     wire start_out_1_34;

     reg [1:0] op_in_1_34;
     wire [1:0] op_out_1_34;

     wire r_1_34;

     reg data_in_1_34;
     wire data_out_1_34;

     reg pivot_in_1_34;
     wire pivot_out_1_34;

     always @(posedge clk) begin
         op_in_1_34 <= op_out_1_33;
         pivot_in_1_34 <= pivot_out_1_33;
         start_in_1_34 <= start_out_1_33;
     end

     always @(posedge clk) begin
         data_in_1_34 <= data_out_0_34;
     end
  
     processor_AB AB_1_34 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_34),
       .start_in   (start_in_1_34),
       .op_in      (op_in_1_34),
       .pivot_in   (pivot_in_1_34),
       .start_out  (start_out_1_34),
       .data_out   (data_out_1_34),
       .op_out     (op_out_1_34),
       .pivot_out  (pivot_out_1_34),
       .r          (r_1_34)
     );

  // row 1, col 35

     reg start_in_1_35;
     wire start_out_1_35;

     reg [1:0] op_in_1_35;
     wire [1:0] op_out_1_35;

     wire r_1_35;

     reg data_in_1_35;
     wire data_out_1_35;

     reg pivot_in_1_35;
     wire pivot_out_1_35;

     always @(posedge clk) begin
         op_in_1_35 <= op_out_1_34;
         pivot_in_1_35 <= pivot_out_1_34;
         start_in_1_35 <= start_out_1_34;
     end

     always @(posedge clk) begin
         data_in_1_35 <= data_out_0_35;
     end
  
     processor_AB AB_1_35 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_35),
       .start_in   (start_in_1_35),
       .op_in      (op_in_1_35),
       .pivot_in   (pivot_in_1_35),
       .start_out  (start_out_1_35),
       .data_out   (data_out_1_35),
       .op_out     (op_out_1_35),
       .pivot_out  (pivot_out_1_35),
       .r          (r_1_35)
     );

  // row 1, col 36

     reg start_in_1_36;
     wire start_out_1_36;

     reg [1:0] op_in_1_36;
     wire [1:0] op_out_1_36;

     wire r_1_36;

     reg data_in_1_36;
     wire data_out_1_36;

     reg pivot_in_1_36;
     wire pivot_out_1_36;

     always @(posedge clk) begin
         op_in_1_36 <= op_out_1_35;
         pivot_in_1_36 <= pivot_out_1_35;
         start_in_1_36 <= start_out_1_35;
     end

     always @(posedge clk) begin
         data_in_1_36 <= data_out_0_36;
     end
  
     processor_AB AB_1_36 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_36),
       .start_in   (start_in_1_36),
       .op_in      (op_in_1_36),
       .pivot_in   (pivot_in_1_36),
       .start_out  (start_out_1_36),
       .data_out   (data_out_1_36),
       .op_out     (op_out_1_36),
       .pivot_out  (pivot_out_1_36),
       .r          (r_1_36)
     );

  // row 1, col 37

     reg start_in_1_37;
     wire start_out_1_37;

     reg [1:0] op_in_1_37;
     wire [1:0] op_out_1_37;

     wire r_1_37;

     reg data_in_1_37;
     wire data_out_1_37;

     reg pivot_in_1_37;
     wire pivot_out_1_37;

     always @(posedge clk) begin
         op_in_1_37 <= op_out_1_36;
         pivot_in_1_37 <= pivot_out_1_36;
         start_in_1_37 <= start_out_1_36;
     end

     always @(posedge clk) begin
         data_in_1_37 <= data_out_0_37;
     end
  
     processor_AB AB_1_37 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_37),
       .start_in   (start_in_1_37),
       .op_in      (op_in_1_37),
       .pivot_in   (pivot_in_1_37),
       .start_out  (start_out_1_37),
       .data_out   (data_out_1_37),
       .op_out     (op_out_1_37),
       .pivot_out  (pivot_out_1_37),
       .r          (r_1_37)
     );

  // row 1, col 38

     reg start_in_1_38;
     wire start_out_1_38;

     reg [1:0] op_in_1_38;
     wire [1:0] op_out_1_38;

     wire r_1_38;

     reg data_in_1_38;
     wire data_out_1_38;

     reg pivot_in_1_38;
     wire pivot_out_1_38;

     always @(posedge clk) begin
         op_in_1_38 <= op_out_1_37;
         pivot_in_1_38 <= pivot_out_1_37;
         start_in_1_38 <= start_out_1_37;
     end

     always @(posedge clk) begin
         data_in_1_38 <= data_out_0_38;
     end
  
     processor_AB AB_1_38 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_38),
       .start_in   (start_in_1_38),
       .op_in      (op_in_1_38),
       .pivot_in   (pivot_in_1_38),
       .start_out  (start_out_1_38),
       .data_out   (data_out_1_38),
       .op_out     (op_out_1_38),
       .pivot_out  (pivot_out_1_38),
       .r          (r_1_38)
     );

  // row 1, col 39

     reg start_in_1_39;
     wire start_out_1_39;

     reg [1:0] op_in_1_39;
     wire [1:0] op_out_1_39;

     wire r_1_39;

     reg data_in_1_39;
     wire data_out_1_39;

     reg pivot_in_1_39;
     wire pivot_out_1_39;

     always @(posedge clk) begin
         op_in_1_39 <= op_out_1_38;
         pivot_in_1_39 <= pivot_out_1_38;
         start_in_1_39 <= start_out_1_38;
     end

     always @(posedge clk) begin
         data_in_1_39 <= data_out_0_39;
     end
  
     processor_AB AB_1_39 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_39),
       .start_in   (start_in_1_39),
       .op_in      (op_in_1_39),
       .pivot_in   (pivot_in_1_39),
       .start_out  (start_out_1_39),
       .data_out   (data_out_1_39),
       .op_out     (op_out_1_39),
       .pivot_out  (pivot_out_1_39),
       .r          (r_1_39)
     );

  // row 1, col 40

     reg start_in_1_40;
     wire start_out_1_40;

     reg [1:0] op_in_1_40;
     wire [1:0] op_out_1_40;

     wire r_1_40;

     reg data_in_1_40;
     wire data_out_1_40;

     reg pivot_in_1_40;
     wire pivot_out_1_40;

     always @(posedge clk) begin
         op_in_1_40 <= op_out_1_39;
         pivot_in_1_40 <= pivot_out_1_39;
         start_in_1_40 <= start_out_1_39;
     end

     always @(posedge clk) begin
         data_in_1_40 <= data_out_0_40;
     end
  
     processor_AB AB_1_40 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_40),
       .start_in   (start_in_1_40),
       .op_in      (op_in_1_40),
       .pivot_in   (pivot_in_1_40),
       .start_out  (start_out_1_40),
       .data_out   (data_out_1_40),
       .op_out     (op_out_1_40),
       .pivot_out  (pivot_out_1_40),
       .r          (r_1_40)
     );

  // row 1, col 41

     reg start_in_1_41;
     wire start_out_1_41;

     reg [1:0] op_in_1_41;
     wire [1:0] op_out_1_41;

     wire r_1_41;

     reg data_in_1_41;
     wire data_out_1_41;

     reg pivot_in_1_41;
     wire pivot_out_1_41;

     always @(posedge clk) begin
         op_in_1_41 <= op_out_1_40;
         pivot_in_1_41 <= pivot_out_1_40;
         start_in_1_41 <= start_out_1_40;
     end

     always @(posedge clk) begin
         data_in_1_41 <= data_out_0_41;
     end
  
     processor_AB AB_1_41 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_41),
       .start_in   (start_in_1_41),
       .op_in      (op_in_1_41),
       .pivot_in   (pivot_in_1_41),
       .start_out  (start_out_1_41),
       .data_out   (data_out_1_41),
       .op_out     (op_out_1_41),
       .pivot_out  (pivot_out_1_41),
       .r          (r_1_41)
     );

  // row 1, col 42

     reg start_in_1_42;
     wire start_out_1_42;

     reg [1:0] op_in_1_42;
     wire [1:0] op_out_1_42;

     wire r_1_42;

     reg data_in_1_42;
     wire data_out_1_42;

     reg pivot_in_1_42;
     wire pivot_out_1_42;

     always @(posedge clk) begin
         op_in_1_42 <= op_out_1_41;
         pivot_in_1_42 <= pivot_out_1_41;
         start_in_1_42 <= start_out_1_41;
     end

     always @(posedge clk) begin
         data_in_1_42 <= data_out_0_42;
     end
  
     processor_AB AB_1_42 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_42),
       .start_in   (start_in_1_42),
       .op_in      (op_in_1_42),
       .pivot_in   (pivot_in_1_42),
       .start_out  (start_out_1_42),
       .data_out   (data_out_1_42),
       .op_out     (op_out_1_42),
       .pivot_out  (pivot_out_1_42),
       .r          (r_1_42)
     );

  // row 1, col 43

     reg start_in_1_43;
     wire start_out_1_43;

     reg [1:0] op_in_1_43;
     wire [1:0] op_out_1_43;

     wire r_1_43;

     reg data_in_1_43;
     wire data_out_1_43;

     reg pivot_in_1_43;
     wire pivot_out_1_43;

     always @(posedge clk) begin
         op_in_1_43 <= op_out_1_42;
         pivot_in_1_43 <= pivot_out_1_42;
         start_in_1_43 <= start_out_1_42;
     end

     always @(posedge clk) begin
         data_in_1_43 <= data_out_0_43;
     end
  
     processor_AB AB_1_43 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_43),
       .start_in   (start_in_1_43),
       .op_in      (op_in_1_43),
       .pivot_in   (pivot_in_1_43),
       .start_out  (start_out_1_43),
       .data_out   (data_out_1_43),
       .op_out     (op_out_1_43),
       .pivot_out  (pivot_out_1_43),
       .r          (r_1_43)
     );

  // row 1, col 44

     reg start_in_1_44;
     wire start_out_1_44;

     reg [1:0] op_in_1_44;
     wire [1:0] op_out_1_44;

     wire r_1_44;

     reg data_in_1_44;
     wire data_out_1_44;

     reg pivot_in_1_44;
     wire pivot_out_1_44;

     always @(posedge clk) begin
         op_in_1_44 <= op_out_1_43;
         pivot_in_1_44 <= pivot_out_1_43;
         start_in_1_44 <= start_out_1_43;
     end

     always @(posedge clk) begin
         data_in_1_44 <= data_out_0_44;
     end
  
     processor_AB AB_1_44 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_44),
       .start_in   (start_in_1_44),
       .op_in      (op_in_1_44),
       .pivot_in   (pivot_in_1_44),
       .start_out  (start_out_1_44),
       .data_out   (data_out_1_44),
       .op_out     (op_out_1_44),
       .pivot_out  (pivot_out_1_44),
       .r          (r_1_44)
     );

  // row 1, col 45

     reg start_in_1_45;
     wire start_out_1_45;

     reg [1:0] op_in_1_45;
     wire [1:0] op_out_1_45;

     wire r_1_45;

     reg data_in_1_45;
     wire data_out_1_45;

     reg pivot_in_1_45;
     wire pivot_out_1_45;

     always @(posedge clk) begin
         op_in_1_45 <= op_out_1_44;
         pivot_in_1_45 <= pivot_out_1_44;
         start_in_1_45 <= start_out_1_44;
     end

     always @(posedge clk) begin
         data_in_1_45 <= data_out_0_45;
     end
  
     processor_AB AB_1_45 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_45),
       .start_in   (start_in_1_45),
       .op_in      (op_in_1_45),
       .pivot_in   (pivot_in_1_45),
       .start_out  (start_out_1_45),
       .data_out   (data_out_1_45),
       .op_out     (op_out_1_45),
       .pivot_out  (pivot_out_1_45),
       .r          (r_1_45)
     );

  // row 1, col 46

     reg start_in_1_46;
     wire start_out_1_46;

     reg [1:0] op_in_1_46;
     wire [1:0] op_out_1_46;

     wire r_1_46;

     reg data_in_1_46;
     wire data_out_1_46;

     reg pivot_in_1_46;
     wire pivot_out_1_46;

     always @(posedge clk) begin
         op_in_1_46 <= op_out_1_45;
         pivot_in_1_46 <= pivot_out_1_45;
         start_in_1_46 <= start_out_1_45;
     end

     always @(posedge clk) begin
         data_in_1_46 <= data_out_0_46;
     end
  
     processor_AB AB_1_46 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_46),
       .start_in   (start_in_1_46),
       .op_in      (op_in_1_46),
       .pivot_in   (pivot_in_1_46),
       .start_out  (start_out_1_46),
       .data_out   (data_out_1_46),
       .op_out     (op_out_1_46),
       .pivot_out  (pivot_out_1_46),
       .r          (r_1_46)
     );

  // row 1, col 47

     reg start_in_1_47;
     wire start_out_1_47;

     reg [1:0] op_in_1_47;
     wire [1:0] op_out_1_47;

     wire r_1_47;

     reg data_in_1_47;
     wire data_out_1_47;

     reg pivot_in_1_47;
     wire pivot_out_1_47;

     always @(posedge clk) begin
         op_in_1_47 <= op_out_1_46;
         pivot_in_1_47 <= pivot_out_1_46;
         start_in_1_47 <= start_out_1_46;
     end

     always @(posedge clk) begin
         data_in_1_47 <= data_out_0_47;
     end
  
     processor_AB AB_1_47 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_47),
       .start_in   (start_in_1_47),
       .op_in      (op_in_1_47),
       .pivot_in   (pivot_in_1_47),
       .start_out  (start_out_1_47),
       .data_out   (data_out_1_47),
       .op_out     (op_out_1_47),
       .pivot_out  (pivot_out_1_47),
       .r          (r_1_47)
     );

  // row 1, col 48

     reg start_in_1_48;
     wire start_out_1_48;

     reg [1:0] op_in_1_48;
     wire [1:0] op_out_1_48;

     wire r_1_48;

     reg data_in_1_48;
     wire data_out_1_48;

     reg pivot_in_1_48;
     wire pivot_out_1_48;

     always @(posedge clk) begin
         op_in_1_48 <= op_out_1_47;
         pivot_in_1_48 <= pivot_out_1_47;
         start_in_1_48 <= start_out_1_47;
     end

     always @(posedge clk) begin
         data_in_1_48 <= data_out_0_48;
     end
  
     processor_AB AB_1_48 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_48),
       .start_in   (start_in_1_48),
       .op_in      (op_in_1_48),
       .pivot_in   (pivot_in_1_48),
       .start_out  (start_out_1_48),
       .data_out   (data_out_1_48),
       .op_out     (op_out_1_48),
       .pivot_out  (pivot_out_1_48),
       .r          (r_1_48)
     );

  // row 1, col 49

     reg start_in_1_49;
     wire start_out_1_49;

     reg [1:0] op_in_1_49;
     wire [1:0] op_out_1_49;

     wire r_1_49;

     reg data_in_1_49;
     wire data_out_1_49;

     reg pivot_in_1_49;
     wire pivot_out_1_49;

     always @(posedge clk) begin
         op_in_1_49 <= op_out_1_48;
         pivot_in_1_49 <= pivot_out_1_48;
         start_in_1_49 <= start_out_1_48;
     end

     always @(posedge clk) begin
         data_in_1_49 <= data_out_0_49;
     end
  
     processor_AB AB_1_49 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_49),
       .start_in   (start_in_1_49),
       .op_in      (op_in_1_49),
       .pivot_in   (pivot_in_1_49),
       .start_out  (start_out_1_49),
       .data_out   (data_out_1_49),
       .op_out     (op_out_1_49),
       .pivot_out  (pivot_out_1_49),
       .r          (r_1_49)
     );

  // row 1, col 50

     reg start_in_1_50;
     wire start_out_1_50;

     reg [1:0] op_in_1_50;
     wire [1:0] op_out_1_50;

     wire r_1_50;

     reg data_in_1_50;
     wire data_out_1_50;

     reg pivot_in_1_50;
     wire pivot_out_1_50;

     always @(posedge clk) begin
         op_in_1_50 <= op_out_1_49;
         pivot_in_1_50 <= pivot_out_1_49;
         start_in_1_50 <= start_out_1_49;
     end

     always @(posedge clk) begin
         data_in_1_50 <= data_out_0_50;
     end
  
     processor_AB AB_1_50 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_50),
       .start_in   (start_in_1_50),
       .op_in      (op_in_1_50),
       .pivot_in   (pivot_in_1_50),
       .start_out  (start_out_1_50),
       .data_out   (data_out_1_50),
       .op_out     (op_out_1_50),
       .pivot_out  (pivot_out_1_50),
       .r          (r_1_50)
     );

  // row 1, col 51

     reg start_in_1_51;
     wire start_out_1_51;

     reg [1:0] op_in_1_51;
     wire [1:0] op_out_1_51;

     wire r_1_51;

     reg data_in_1_51;
     wire data_out_1_51;

     reg pivot_in_1_51;
     wire pivot_out_1_51;

     always @(posedge clk) begin
         op_in_1_51 <= op_out_1_50;
         pivot_in_1_51 <= pivot_out_1_50;
         start_in_1_51 <= start_out_1_50;
     end

     always @(posedge clk) begin
         data_in_1_51 <= data_out_0_51;
     end
  
     processor_AB AB_1_51 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_51),
       .start_in   (start_in_1_51),
       .op_in      (op_in_1_51),
       .pivot_in   (pivot_in_1_51),
       .start_out  (start_out_1_51),
       .data_out   (data_out_1_51),
       .op_out     (op_out_1_51),
       .pivot_out  (pivot_out_1_51),
       .r          (r_1_51)
     );

  // row 1, col 52

     reg start_in_1_52;
     wire start_out_1_52;

     reg [1:0] op_in_1_52;
     wire [1:0] op_out_1_52;

     wire r_1_52;

     reg data_in_1_52;
     wire data_out_1_52;

     reg pivot_in_1_52;
     wire pivot_out_1_52;

     always @(posedge clk) begin
         op_in_1_52 <= op_out_1_51;
         pivot_in_1_52 <= pivot_out_1_51;
         start_in_1_52 <= start_out_1_51;
     end

     always @(posedge clk) begin
         data_in_1_52 <= data_out_0_52;
     end
  
     processor_AB AB_1_52 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_52),
       .start_in   (start_in_1_52),
       .op_in      (op_in_1_52),
       .pivot_in   (pivot_in_1_52),
       .start_out  (start_out_1_52),
       .data_out   (data_out_1_52),
       .op_out     (op_out_1_52),
       .pivot_out  (pivot_out_1_52),
       .r          (r_1_52)
     );

  // row 1, col 53

     reg start_in_1_53;
     wire start_out_1_53;

     reg [1:0] op_in_1_53;
     wire [1:0] op_out_1_53;

     wire r_1_53;

     reg data_in_1_53;
     wire data_out_1_53;

     reg pivot_in_1_53;
     wire pivot_out_1_53;

     always @(posedge clk) begin
         op_in_1_53 <= op_out_1_52;
         pivot_in_1_53 <= pivot_out_1_52;
         start_in_1_53 <= start_out_1_52;
     end

     always @(posedge clk) begin
         data_in_1_53 <= data_out_0_53;
     end
  
     processor_AB AB_1_53 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_53),
       .start_in   (start_in_1_53),
       .op_in      (op_in_1_53),
       .pivot_in   (pivot_in_1_53),
       .start_out  (start_out_1_53),
       .data_out   (data_out_1_53),
       .op_out     (op_out_1_53),
       .pivot_out  (pivot_out_1_53),
       .r          (r_1_53)
     );

  // row 1, col 54

     reg start_in_1_54;
     wire start_out_1_54;

     reg [1:0] op_in_1_54;
     wire [1:0] op_out_1_54;

     wire r_1_54;

     reg data_in_1_54;
     wire data_out_1_54;

     reg pivot_in_1_54;
     wire pivot_out_1_54;

     always @(posedge clk) begin
         op_in_1_54 <= op_out_1_53;
         pivot_in_1_54 <= pivot_out_1_53;
         start_in_1_54 <= start_out_1_53;
     end

     always @(posedge clk) begin
         data_in_1_54 <= data_out_0_54;
     end
  
     processor_AB AB_1_54 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_54),
       .start_in   (start_in_1_54),
       .op_in      (op_in_1_54),
       .pivot_in   (pivot_in_1_54),
       .start_out  (start_out_1_54),
       .data_out   (data_out_1_54),
       .op_out     (op_out_1_54),
       .pivot_out  (pivot_out_1_54),
       .r          (r_1_54)
     );

  // row 1, col 55

     reg start_in_1_55;
     wire start_out_1_55;

     reg [1:0] op_in_1_55;
     wire [1:0] op_out_1_55;

     wire r_1_55;

     reg data_in_1_55;
     wire data_out_1_55;

     reg pivot_in_1_55;
     wire pivot_out_1_55;

     always @(posedge clk) begin
         op_in_1_55 <= op_out_1_54;
         pivot_in_1_55 <= pivot_out_1_54;
         start_in_1_55 <= start_out_1_54;
     end

     always @(posedge clk) begin
         data_in_1_55 <= data_out_0_55;
     end
  
     processor_AB AB_1_55 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_55),
       .start_in   (start_in_1_55),
       .op_in      (op_in_1_55),
       .pivot_in   (pivot_in_1_55),
       .start_out  (start_out_1_55),
       .data_out   (data_out_1_55),
       .op_out     (op_out_1_55),
       .pivot_out  (pivot_out_1_55),
       .r          (r_1_55)
     );

  // row 1, col 56

     reg start_in_1_56;
     wire start_out_1_56;

     reg [1:0] op_in_1_56;
     wire [1:0] op_out_1_56;

     wire r_1_56;

     reg data_in_1_56;
     wire data_out_1_56;

     reg pivot_in_1_56;
     wire pivot_out_1_56;

     always @(posedge clk) begin
         op_in_1_56 <= op_out_1_55;
         pivot_in_1_56 <= pivot_out_1_55;
         start_in_1_56 <= start_out_1_55;
     end

     always @(posedge clk) begin
         data_in_1_56 <= data_out_0_56;
     end
  
     processor_AB AB_1_56 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_56),
       .start_in   (start_in_1_56),
       .op_in      (op_in_1_56),
       .pivot_in   (pivot_in_1_56),
       .start_out  (start_out_1_56),
       .data_out   (data_out_1_56),
       .op_out     (op_out_1_56),
       .pivot_out  (pivot_out_1_56),
       .r          (r_1_56)
     );

  // row 1, col 57

     reg start_in_1_57;
     wire start_out_1_57;

     reg [1:0] op_in_1_57;
     wire [1:0] op_out_1_57;

     wire r_1_57;

     reg data_in_1_57;
     wire data_out_1_57;

     reg pivot_in_1_57;
     wire pivot_out_1_57;

     always @(posedge clk) begin
         op_in_1_57 <= op_out_1_56;
         pivot_in_1_57 <= pivot_out_1_56;
         start_in_1_57 <= start_out_1_56;
     end

     always @(posedge clk) begin
         data_in_1_57 <= data_out_0_57;
     end
  
     processor_AB AB_1_57 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_57),
       .start_in   (start_in_1_57),
       .op_in      (op_in_1_57),
       .pivot_in   (pivot_in_1_57),
       .start_out  (start_out_1_57),
       .data_out   (data_out_1_57),
       .op_out     (op_out_1_57),
       .pivot_out  (pivot_out_1_57),
       .r          (r_1_57)
     );

  // row 1, col 58

     reg start_in_1_58;
     wire start_out_1_58;

     reg [1:0] op_in_1_58;
     wire [1:0] op_out_1_58;

     wire r_1_58;

     reg data_in_1_58;
     wire data_out_1_58;

     reg pivot_in_1_58;
     wire pivot_out_1_58;

     always @(posedge clk) begin
         op_in_1_58 <= op_out_1_57;
         pivot_in_1_58 <= pivot_out_1_57;
         start_in_1_58 <= start_out_1_57;
     end

     always @(posedge clk) begin
         data_in_1_58 <= data_out_0_58;
     end
  
     processor_AB AB_1_58 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_58),
       .start_in   (start_in_1_58),
       .op_in      (op_in_1_58),
       .pivot_in   (pivot_in_1_58),
       .start_out  (start_out_1_58),
       .data_out   (data_out_1_58),
       .op_out     (op_out_1_58),
       .pivot_out  (pivot_out_1_58),
       .r          (r_1_58)
     );

  // row 1, col 59

     reg start_in_1_59;
     wire start_out_1_59;

     reg [1:0] op_in_1_59;
     wire [1:0] op_out_1_59;

     wire r_1_59;

     reg data_in_1_59;
     wire data_out_1_59;

     reg pivot_in_1_59;
     wire pivot_out_1_59;

     always @(posedge clk) begin
         op_in_1_59 <= op_out_1_58;
         pivot_in_1_59 <= pivot_out_1_58;
         start_in_1_59 <= start_out_1_58;
     end

     always @(posedge clk) begin
         data_in_1_59 <= data_out_0_59;
     end
  
     processor_AB AB_1_59 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_59),
       .start_in   (start_in_1_59),
       .op_in      (op_in_1_59),
       .pivot_in   (pivot_in_1_59),
       .start_out  (start_out_1_59),
       .data_out   (data_out_1_59),
       .op_out     (op_out_1_59),
       .pivot_out  (pivot_out_1_59),
       .r          (r_1_59)
     );

  // row 1, col 60

     reg start_in_1_60;
     wire start_out_1_60;

     reg [1:0] op_in_1_60;
     wire [1:0] op_out_1_60;

     wire r_1_60;

     reg data_in_1_60;
     wire data_out_1_60;

     reg pivot_in_1_60;
     wire pivot_out_1_60;

     always @(posedge clk) begin
         op_in_1_60 <= op_out_1_59;
         pivot_in_1_60 <= pivot_out_1_59;
         start_in_1_60 <= start_out_1_59;
     end

     always @(posedge clk) begin
         data_in_1_60 <= data_out_0_60;
     end
  
     processor_AB AB_1_60 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_60),
       .start_in   (start_in_1_60),
       .op_in      (op_in_1_60),
       .pivot_in   (pivot_in_1_60),
       .start_out  (start_out_1_60),
       .data_out   (data_out_1_60),
       .op_out     (op_out_1_60),
       .pivot_out  (pivot_out_1_60),
       .r          (r_1_60)
     );

  // row 1, col 61

     reg start_in_1_61;
     wire start_out_1_61;

     reg [1:0] op_in_1_61;
     wire [1:0] op_out_1_61;

     wire r_1_61;

     reg data_in_1_61;
     wire data_out_1_61;

     reg pivot_in_1_61;
     wire pivot_out_1_61;

     always @(posedge clk) begin
         op_in_1_61 <= op_out_1_60;
         pivot_in_1_61 <= pivot_out_1_60;
         start_in_1_61 <= start_out_1_60;
     end

     always @(posedge clk) begin
         data_in_1_61 <= data_out_0_61;
     end
  
     processor_AB AB_1_61 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_61),
       .start_in   (start_in_1_61),
       .op_in      (op_in_1_61),
       .pivot_in   (pivot_in_1_61),
       .start_out  (start_out_1_61),
       .data_out   (data_out_1_61),
       .op_out     (op_out_1_61),
       .pivot_out  (pivot_out_1_61),
       .r          (r_1_61)
     );

  // row 1, col 62

     reg start_in_1_62;
     wire start_out_1_62;

     reg [1:0] op_in_1_62;
     wire [1:0] op_out_1_62;

     wire r_1_62;

     reg data_in_1_62;
     wire data_out_1_62;

     reg pivot_in_1_62;
     wire pivot_out_1_62;

     always @(posedge clk) begin
         op_in_1_62 <= op_out_1_61;
         pivot_in_1_62 <= pivot_out_1_61;
         start_in_1_62 <= start_out_1_61;
     end

     always @(posedge clk) begin
         data_in_1_62 <= data_out_0_62;
     end
  
     processor_AB AB_1_62 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_62),
       .start_in   (start_in_1_62),
       .op_in      (op_in_1_62),
       .pivot_in   (pivot_in_1_62),
       .start_out  (start_out_1_62),
       .data_out   (data_out_1_62),
       .op_out     (op_out_1_62),
       .pivot_out  (pivot_out_1_62),
       .r          (r_1_62)
     );

  // row 1, col 63

     reg start_in_1_63;
     wire start_out_1_63;

     reg [1:0] op_in_1_63;
     wire [1:0] op_out_1_63;

     wire r_1_63;

     reg data_in_1_63;
     wire data_out_1_63;

     reg pivot_in_1_63;
     wire pivot_out_1_63;

     always @(posedge clk) begin
         op_in_1_63 <= op_out_1_62;
         pivot_in_1_63 <= pivot_out_1_62;
         start_in_1_63 <= start_out_1_62;
     end

     always @(posedge clk) begin
         data_in_1_63 <= data_out_0_63;
     end
  
     processor_AB AB_1_63 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_63),
       .start_in   (start_in_1_63),
       .op_in      (op_in_1_63),
       .pivot_in   (pivot_in_1_63),
       .start_out  (start_out_1_63),
       .data_out   (data_out_1_63),
       .op_out     (op_out_1_63),
       .pivot_out  (pivot_out_1_63),
       .r          (r_1_63)
     );

  // row 1, col 64

     reg start_in_1_64;
     wire start_out_1_64;

     reg [1:0] op_in_1_64;
     wire [1:0] op_out_1_64;

     wire r_1_64;

     reg data_in_1_64;
     wire data_out_1_64;

     reg pivot_in_1_64;
     wire pivot_out_1_64;

     always @(posedge clk) begin
         op_in_1_64 <= op_out_1_63;
         pivot_in_1_64 <= pivot_out_1_63;
         start_in_1_64 <= start_out_1_63;
     end

     always @(posedge clk) begin
         data_in_1_64 <= data_out_0_64;
     end
  
     processor_AB AB_1_64 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_64),
       .start_in   (start_in_1_64),
       .op_in      (op_in_1_64),
       .pivot_in   (pivot_in_1_64),
       .start_out  (start_out_1_64),
       .data_out   (data_out_1_64),
       .op_out     (op_out_1_64),
       .pivot_out  (pivot_out_1_64),
       .r          (r_1_64)
     );

  // row 1, col 65

     reg start_in_1_65;
     wire start_out_1_65;

     reg [1:0] op_in_1_65;
     wire [1:0] op_out_1_65;

     wire r_1_65;

     reg data_in_1_65;
     wire data_out_1_65;

     reg pivot_in_1_65;
     wire pivot_out_1_65;

     always @(posedge clk) begin
         op_in_1_65 <= op_out_1_64;
         pivot_in_1_65 <= pivot_out_1_64;
         start_in_1_65 <= start_out_1_64;
     end

     always @(posedge clk) begin
         data_in_1_65 <= data_out_0_65;
     end
  
     processor_AB AB_1_65 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_65),
       .start_in   (start_in_1_65),
       .op_in      (op_in_1_65),
       .pivot_in   (pivot_in_1_65),
       .start_out  (start_out_1_65),
       .data_out   (data_out_1_65),
       .op_out     (op_out_1_65),
       .pivot_out  (pivot_out_1_65),
       .r          (r_1_65)
     );

  // row 1, col 66

     reg start_in_1_66;
     wire start_out_1_66;

     reg [1:0] op_in_1_66;
     wire [1:0] op_out_1_66;

     wire r_1_66;

     reg data_in_1_66;
     wire data_out_1_66;

     reg pivot_in_1_66;
     wire pivot_out_1_66;

     always @(posedge clk) begin
         op_in_1_66 <= op_out_1_65;
         pivot_in_1_66 <= pivot_out_1_65;
         start_in_1_66 <= start_out_1_65;
     end

     always @(posedge clk) begin
         data_in_1_66 <= data_out_0_66;
     end
  
     processor_AB AB_1_66 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_66),
       .start_in   (start_in_1_66),
       .op_in      (op_in_1_66),
       .pivot_in   (pivot_in_1_66),
       .start_out  (start_out_1_66),
       .data_out   (data_out_1_66),
       .op_out     (op_out_1_66),
       .pivot_out  (pivot_out_1_66),
       .r          (r_1_66)
     );

  // row 1, col 67

     reg start_in_1_67;
     wire start_out_1_67;

     reg [1:0] op_in_1_67;
     wire [1:0] op_out_1_67;

     wire r_1_67;

     reg data_in_1_67;
     wire data_out_1_67;

     reg pivot_in_1_67;
     wire pivot_out_1_67;

     always @(posedge clk) begin
         op_in_1_67 <= op_out_1_66;
         pivot_in_1_67 <= pivot_out_1_66;
         start_in_1_67 <= start_out_1_66;
     end

     always @(posedge clk) begin
         data_in_1_67 <= data_out_0_67;
     end
  
     processor_AB AB_1_67 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_67),
       .start_in   (start_in_1_67),
       .op_in      (op_in_1_67),
       .pivot_in   (pivot_in_1_67),
       .start_out  (start_out_1_67),
       .data_out   (data_out_1_67),
       .op_out     (op_out_1_67),
       .pivot_out  (pivot_out_1_67),
       .r          (r_1_67)
     );

  // row 1, col 68

     reg start_in_1_68;
     wire start_out_1_68;

     reg [1:0] op_in_1_68;
     wire [1:0] op_out_1_68;

     wire r_1_68;

     reg data_in_1_68;
     wire data_out_1_68;

     reg pivot_in_1_68;
     wire pivot_out_1_68;

     always @(posedge clk) begin
         op_in_1_68 <= op_out_1_67;
         pivot_in_1_68 <= pivot_out_1_67;
         start_in_1_68 <= start_out_1_67;
     end

     always @(posedge clk) begin
         data_in_1_68 <= data_out_0_68;
     end
  
     processor_AB AB_1_68 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_68),
       .start_in   (start_in_1_68),
       .op_in      (op_in_1_68),
       .pivot_in   (pivot_in_1_68),
       .start_out  (start_out_1_68),
       .data_out   (data_out_1_68),
       .op_out     (op_out_1_68),
       .pivot_out  (pivot_out_1_68),
       .r          (r_1_68)
     );

  // row 1, col 69

     reg start_in_1_69;
     wire start_out_1_69;

     reg [1:0] op_in_1_69;
     wire [1:0] op_out_1_69;

     wire r_1_69;

     reg data_in_1_69;
     wire data_out_1_69;

     reg pivot_in_1_69;
     wire pivot_out_1_69;

     always @(posedge clk) begin
         op_in_1_69 <= op_out_1_68;
         pivot_in_1_69 <= pivot_out_1_68;
         start_in_1_69 <= start_out_1_68;
     end

     always @(posedge clk) begin
         data_in_1_69 <= data_out_0_69;
     end
  
     processor_AB AB_1_69 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_69),
       .start_in   (start_in_1_69),
       .op_in      (op_in_1_69),
       .pivot_in   (pivot_in_1_69),
       .start_out  (start_out_1_69),
       .data_out   (data_out_1_69),
       .op_out     (op_out_1_69),
       .pivot_out  (pivot_out_1_69),
       .r          (r_1_69)
     );

  // row 1, col 70

     reg start_in_1_70;
     wire start_out_1_70;

     reg [1:0] op_in_1_70;
     wire [1:0] op_out_1_70;

     wire r_1_70;

     reg data_in_1_70;
     wire data_out_1_70;

     reg pivot_in_1_70;
     wire pivot_out_1_70;

     always @(posedge clk) begin
         op_in_1_70 <= op_out_1_69;
         pivot_in_1_70 <= pivot_out_1_69;
         start_in_1_70 <= start_out_1_69;
     end

     always @(posedge clk) begin
         data_in_1_70 <= data_out_0_70;
     end
  
     processor_AB AB_1_70 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_70),
       .start_in   (start_in_1_70),
       .op_in      (op_in_1_70),
       .pivot_in   (pivot_in_1_70),
       .start_out  (start_out_1_70),
       .data_out   (data_out_1_70),
       .op_out     (op_out_1_70),
       .pivot_out  (pivot_out_1_70),
       .r          (r_1_70)
     );

  // row 1, col 71

     reg start_in_1_71;
     wire start_out_1_71;

     reg [1:0] op_in_1_71;
     wire [1:0] op_out_1_71;

     wire r_1_71;

     reg data_in_1_71;
     wire data_out_1_71;

     reg pivot_in_1_71;
     wire pivot_out_1_71;

     always @(posedge clk) begin
         op_in_1_71 <= op_out_1_70;
         pivot_in_1_71 <= pivot_out_1_70;
         start_in_1_71 <= start_out_1_70;
     end

     always @(posedge clk) begin
         data_in_1_71 <= data_out_0_71;
     end
  
     processor_AB AB_1_71 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_71),
       .start_in   (start_in_1_71),
       .op_in      (op_in_1_71),
       .pivot_in   (pivot_in_1_71),
       .start_out  (start_out_1_71),
       .data_out   (data_out_1_71),
       .op_out     (op_out_1_71),
       .pivot_out  (pivot_out_1_71),
       .r          (r_1_71)
     );

  // row 1, col 72

     reg start_in_1_72;
     wire start_out_1_72;

     reg [1:0] op_in_1_72;
     wire [1:0] op_out_1_72;

     wire r_1_72;

     reg data_in_1_72;
     wire data_out_1_72;

     reg pivot_in_1_72;
     wire pivot_out_1_72;

     always @(posedge clk) begin
         op_in_1_72 <= op_out_1_71;
         pivot_in_1_72 <= pivot_out_1_71;
         start_in_1_72 <= start_out_1_71;
     end

     always @(posedge clk) begin
         data_in_1_72 <= data_out_0_72;
     end
  
     processor_AB AB_1_72 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_72),
       .start_in   (start_in_1_72),
       .op_in      (op_in_1_72),
       .pivot_in   (pivot_in_1_72),
       .start_out  (start_out_1_72),
       .data_out   (data_out_1_72),
       .op_out     (op_out_1_72),
       .pivot_out  (pivot_out_1_72),
       .r          (r_1_72)
     );

  // row 1, col 73

     reg start_in_1_73;
     wire start_out_1_73;

     reg [1:0] op_in_1_73;
     wire [1:0] op_out_1_73;

     wire r_1_73;

     reg data_in_1_73;
     wire data_out_1_73;

     reg pivot_in_1_73;
     wire pivot_out_1_73;

     always @(posedge clk) begin
         op_in_1_73 <= op_out_1_72;
         pivot_in_1_73 <= pivot_out_1_72;
         start_in_1_73 <= start_out_1_72;
     end

     always @(posedge clk) begin
         data_in_1_73 <= data_out_0_73;
     end
  
     processor_AB AB_1_73 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_73),
       .start_in   (start_in_1_73),
       .op_in      (op_in_1_73),
       .pivot_in   (pivot_in_1_73),
       .start_out  (start_out_1_73),
       .data_out   (data_out_1_73),
       .op_out     (op_out_1_73),
       .pivot_out  (pivot_out_1_73),
       .r          (r_1_73)
     );

  // row 1, col 74

     reg start_in_1_74;
     wire start_out_1_74;

     reg [1:0] op_in_1_74;
     wire [1:0] op_out_1_74;

     wire r_1_74;

     reg data_in_1_74;
     wire data_out_1_74;

     reg pivot_in_1_74;
     wire pivot_out_1_74;

     always @(posedge clk) begin
         op_in_1_74 <= op_out_1_73;
         pivot_in_1_74 <= pivot_out_1_73;
         start_in_1_74 <= start_out_1_73;
     end

     always @(posedge clk) begin
         data_in_1_74 <= data_out_0_74;
     end
  
     processor_AB AB_1_74 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_74),
       .start_in   (start_in_1_74),
       .op_in      (op_in_1_74),
       .pivot_in   (pivot_in_1_74),
       .start_out  (start_out_1_74),
       .data_out   (data_out_1_74),
       .op_out     (op_out_1_74),
       .pivot_out  (pivot_out_1_74),
       .r          (r_1_74)
     );

  // row 1, col 75

     reg start_in_1_75;
     wire start_out_1_75;

     reg [1:0] op_in_1_75;
     wire [1:0] op_out_1_75;

     wire r_1_75;

     reg data_in_1_75;
     wire data_out_1_75;

     reg pivot_in_1_75;
     wire pivot_out_1_75;

     always @(posedge clk) begin
         op_in_1_75 <= op_out_1_74;
         pivot_in_1_75 <= pivot_out_1_74;
         start_in_1_75 <= start_out_1_74;
     end

     always @(posedge clk) begin
         data_in_1_75 <= data_out_0_75;
     end
  
     processor_AB AB_1_75 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_75),
       .start_in   (start_in_1_75),
       .op_in      (op_in_1_75),
       .pivot_in   (pivot_in_1_75),
       .start_out  (start_out_1_75),
       .data_out   (data_out_1_75),
       .op_out     (op_out_1_75),
       .pivot_out  (pivot_out_1_75),
       .r          (r_1_75)
     );

  // row 1, col 76

     reg start_in_1_76;
     wire start_out_1_76;

     reg [1:0] op_in_1_76;
     wire [1:0] op_out_1_76;

     wire r_1_76;

     reg data_in_1_76;
     wire data_out_1_76;

     reg pivot_in_1_76;
     wire pivot_out_1_76;

     always @(posedge clk) begin
         op_in_1_76 <= op_out_1_75;
         pivot_in_1_76 <= pivot_out_1_75;
         start_in_1_76 <= start_out_1_75;
     end

     always @(posedge clk) begin
         data_in_1_76 <= data_out_0_76;
     end
  
     processor_AB AB_1_76 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_76),
       .start_in   (start_in_1_76),
       .op_in      (op_in_1_76),
       .pivot_in   (pivot_in_1_76),
       .start_out  (start_out_1_76),
       .data_out   (data_out_1_76),
       .op_out     (op_out_1_76),
       .pivot_out  (pivot_out_1_76),
       .r          (r_1_76)
     );

  // row 1, col 77

     reg start_in_1_77;
     wire start_out_1_77;

     reg [1:0] op_in_1_77;
     wire [1:0] op_out_1_77;

     wire r_1_77;

     reg data_in_1_77;
     wire data_out_1_77;

     reg pivot_in_1_77;
     wire pivot_out_1_77;

     always @(posedge clk) begin
         op_in_1_77 <= op_out_1_76;
         pivot_in_1_77 <= pivot_out_1_76;
         start_in_1_77 <= start_out_1_76;
     end

     always @(posedge clk) begin
         data_in_1_77 <= data_out_0_77;
     end
  
     processor_AB AB_1_77 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_77),
       .start_in   (start_in_1_77),
       .op_in      (op_in_1_77),
       .pivot_in   (pivot_in_1_77),
       .start_out  (start_out_1_77),
       .data_out   (data_out_1_77),
       .op_out     (op_out_1_77),
       .pivot_out  (pivot_out_1_77),
       .r          (r_1_77)
     );

  // row 1, col 78

     reg start_in_1_78;
     wire start_out_1_78;

     reg [1:0] op_in_1_78;
     wire [1:0] op_out_1_78;

     wire r_1_78;

     reg data_in_1_78;
     wire data_out_1_78;

     reg pivot_in_1_78;
     wire pivot_out_1_78;

     always @(posedge clk) begin
         op_in_1_78 <= op_out_1_77;
         pivot_in_1_78 <= pivot_out_1_77;
         start_in_1_78 <= start_out_1_77;
     end

     always @(posedge clk) begin
         data_in_1_78 <= data_out_0_78;
     end
  
     processor_AB AB_1_78 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_78),
       .start_in   (start_in_1_78),
       .op_in      (op_in_1_78),
       .pivot_in   (pivot_in_1_78),
       .start_out  (start_out_1_78),
       .data_out   (data_out_1_78),
       .op_out     (op_out_1_78),
       .pivot_out  (pivot_out_1_78),
       .r          (r_1_78)
     );

  // row 1, col 79

     reg start_in_1_79;
     wire start_out_1_79;

     reg [1:0] op_in_1_79;
     wire [1:0] op_out_1_79;

     wire r_1_79;

     reg data_in_1_79;
     wire data_out_1_79;

     reg pivot_in_1_79;
     wire pivot_out_1_79;

     always @(posedge clk) begin
         op_in_1_79 <= op_out_1_78;
         pivot_in_1_79 <= pivot_out_1_78;
         start_in_1_79 <= start_out_1_78;
     end

     always @(posedge clk) begin
         data_in_1_79 <= data_out_0_79;
     end
  
     processor_AB AB_1_79 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_79),
       .start_in   (start_in_1_79),
       .op_in      (op_in_1_79),
       .pivot_in   (pivot_in_1_79),
       .start_out  (start_out_1_79),
       .data_out   (data_out_1_79),
       .op_out     (op_out_1_79),
       .pivot_out  (pivot_out_1_79),
       .r          (r_1_79)
     );

  // row 1, col 80

     reg start_in_1_80;
     wire start_out_1_80;

     reg [1:0] op_in_1_80;
     wire [1:0] op_out_1_80;

     wire r_1_80;

     reg data_in_1_80;
     wire data_out_1_80;

     reg pivot_in_1_80;
     wire pivot_out_1_80;

     always @(posedge clk) begin
         op_in_1_80 <= op_out_1_79;
         pivot_in_1_80 <= pivot_out_1_79;
         start_in_1_80 <= start_out_1_79;
     end

     always @(posedge clk) begin
         data_in_1_80 <= data_out_0_80;
     end
  
     processor_AB AB_1_80 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_80),
       .start_in   (start_in_1_80),
       .op_in      (op_in_1_80),
       .pivot_in   (pivot_in_1_80),
       .start_out  (start_out_1_80),
       .data_out   (data_out_1_80),
       .op_out     (op_out_1_80),
       .pivot_out  (pivot_out_1_80),
       .r          (r_1_80)
     );

  // row 1, col 81

     reg start_in_1_81;
     wire start_out_1_81;

     reg [1:0] op_in_1_81;
     wire [1:0] op_out_1_81;

     wire r_1_81;

     reg data_in_1_81;
     wire data_out_1_81;

     reg pivot_in_1_81;
     wire pivot_out_1_81;

     always @(posedge clk) begin
         op_in_1_81 <= op_out_1_80;
         pivot_in_1_81 <= pivot_out_1_80;
         start_in_1_81 <= start_out_1_80;
     end

     always @(posedge clk) begin
         data_in_1_81 <= data_out_0_81;
     end
  
     processor_AB AB_1_81 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_81),
       .start_in   (start_in_1_81),
       .op_in      (op_in_1_81),
       .pivot_in   (pivot_in_1_81),
       .start_out  (start_out_1_81),
       .data_out   (data_out_1_81),
       .op_out     (op_out_1_81),
       .pivot_out  (pivot_out_1_81),
       .r          (r_1_81)
     );

  // row 1, col 82

     reg start_in_1_82;
     wire start_out_1_82;

     reg [1:0] op_in_1_82;
     wire [1:0] op_out_1_82;

     wire r_1_82;

     reg data_in_1_82;
     wire data_out_1_82;

     reg pivot_in_1_82;
     wire pivot_out_1_82;

     always @(posedge clk) begin
         op_in_1_82 <= op_out_1_81;
         pivot_in_1_82 <= pivot_out_1_81;
         start_in_1_82 <= start_out_1_81;
     end

     always @(posedge clk) begin
         data_in_1_82 <= data_out_0_82;
     end
  
     processor_AB AB_1_82 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_82),
       .start_in   (start_in_1_82),
       .op_in      (op_in_1_82),
       .pivot_in   (pivot_in_1_82),
       .start_out  (start_out_1_82),
       .data_out   (data_out_1_82),
       .op_out     (op_out_1_82),
       .pivot_out  (pivot_out_1_82),
       .r          (r_1_82)
     );

  // row 1, col 83

     reg start_in_1_83;
     wire start_out_1_83;

     reg [1:0] op_in_1_83;
     wire [1:0] op_out_1_83;

     wire r_1_83;

     reg data_in_1_83;
     wire data_out_1_83;

     reg pivot_in_1_83;
     wire pivot_out_1_83;

     always @(posedge clk) begin
         op_in_1_83 <= op_out_1_82;
         pivot_in_1_83 <= pivot_out_1_82;
         start_in_1_83 <= start_out_1_82;
     end

     always @(posedge clk) begin
         data_in_1_83 <= data_out_0_83;
     end
  
     processor_AB AB_1_83 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_83),
       .start_in   (start_in_1_83),
       .op_in      (op_in_1_83),
       .pivot_in   (pivot_in_1_83),
       .start_out  (start_out_1_83),
       .data_out   (data_out_1_83),
       .op_out     (op_out_1_83),
       .pivot_out  (pivot_out_1_83),
       .r          (r_1_83)
     );

  // row 1, col 84

     reg start_in_1_84;
     wire start_out_1_84;

     reg [1:0] op_in_1_84;
     wire [1:0] op_out_1_84;

     wire r_1_84;

     reg data_in_1_84;
     wire data_out_1_84;

     reg pivot_in_1_84;
     wire pivot_out_1_84;

     always @(posedge clk) begin
         op_in_1_84 <= op_out_1_83;
         pivot_in_1_84 <= pivot_out_1_83;
         start_in_1_84 <= start_out_1_83;
     end

     always @(posedge clk) begin
         data_in_1_84 <= data_out_0_84;
     end
  
     processor_AB AB_1_84 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_84),
       .start_in   (start_in_1_84),
       .op_in      (op_in_1_84),
       .pivot_in   (pivot_in_1_84),
       .start_out  (start_out_1_84),
       .data_out   (data_out_1_84),
       .op_out     (op_out_1_84),
       .pivot_out  (pivot_out_1_84),
       .r          (r_1_84)
     );

  // row 1, col 85

     reg start_in_1_85;
     wire start_out_1_85;

     reg [1:0] op_in_1_85;
     wire [1:0] op_out_1_85;

     wire r_1_85;

     reg data_in_1_85;
     wire data_out_1_85;

     reg pivot_in_1_85;
     wire pivot_out_1_85;

     always @(posedge clk) begin
         op_in_1_85 <= op_out_1_84;
         pivot_in_1_85 <= pivot_out_1_84;
         start_in_1_85 <= start_out_1_84;
     end

     always @(posedge clk) begin
         data_in_1_85 <= data_out_0_85;
     end
  
     processor_AB AB_1_85 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_85),
       .start_in   (start_in_1_85),
       .op_in      (op_in_1_85),
       .pivot_in   (pivot_in_1_85),
       .start_out  (start_out_1_85),
       .data_out   (data_out_1_85),
       .op_out     (op_out_1_85),
       .pivot_out  (pivot_out_1_85),
       .r          (r_1_85)
     );

  // row 1, col 86

     reg start_in_1_86;
     wire start_out_1_86;

     reg [1:0] op_in_1_86;
     wire [1:0] op_out_1_86;

     wire r_1_86;

     reg data_in_1_86;
     wire data_out_1_86;

     reg pivot_in_1_86;
     wire pivot_out_1_86;

     always @(posedge clk) begin
         op_in_1_86 <= op_out_1_85;
         pivot_in_1_86 <= pivot_out_1_85;
         start_in_1_86 <= start_out_1_85;
     end

     always @(posedge clk) begin
         data_in_1_86 <= data_out_0_86;
     end
  
     processor_AB AB_1_86 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_86),
       .start_in   (start_in_1_86),
       .op_in      (op_in_1_86),
       .pivot_in   (pivot_in_1_86),
       .start_out  (start_out_1_86),
       .data_out   (data_out_1_86),
       .op_out     (op_out_1_86),
       .pivot_out  (pivot_out_1_86),
       .r          (r_1_86)
     );

  // row 1, col 87

     reg start_in_1_87;
     wire start_out_1_87;

     reg [1:0] op_in_1_87;
     wire [1:0] op_out_1_87;

     wire r_1_87;

     reg data_in_1_87;
     wire data_out_1_87;

     reg pivot_in_1_87;
     wire pivot_out_1_87;

     always @(posedge clk) begin
         op_in_1_87 <= op_out_1_86;
         pivot_in_1_87 <= pivot_out_1_86;
         start_in_1_87 <= start_out_1_86;
     end

     always @(posedge clk) begin
         data_in_1_87 <= data_out_0_87;
     end
  
     processor_AB AB_1_87 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_87),
       .start_in   (start_in_1_87),
       .op_in      (op_in_1_87),
       .pivot_in   (pivot_in_1_87),
       .start_out  (start_out_1_87),
       .data_out   (data_out_1_87),
       .op_out     (op_out_1_87),
       .pivot_out  (pivot_out_1_87),
       .r          (r_1_87)
     );

  // row 1, col 88

     reg start_in_1_88;
     wire start_out_1_88;

     reg [1:0] op_in_1_88;
     wire [1:0] op_out_1_88;

     wire r_1_88;

     reg data_in_1_88;
     wire data_out_1_88;

     reg pivot_in_1_88;
     wire pivot_out_1_88;

     always @(posedge clk) begin
         op_in_1_88 <= op_out_1_87;
         pivot_in_1_88 <= pivot_out_1_87;
         start_in_1_88 <= start_out_1_87;
     end

     always @(posedge clk) begin
         data_in_1_88 <= data_out_0_88;
     end
  
     processor_AB AB_1_88 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_88),
       .start_in   (start_in_1_88),
       .op_in      (op_in_1_88),
       .pivot_in   (pivot_in_1_88),
       .start_out  (start_out_1_88),
       .data_out   (data_out_1_88),
       .op_out     (op_out_1_88),
       .pivot_out  (pivot_out_1_88),
       .r          (r_1_88)
     );

  // row 1, col 89

     reg start_in_1_89;
     wire start_out_1_89;

     reg [1:0] op_in_1_89;
     wire [1:0] op_out_1_89;

     wire r_1_89;

     reg data_in_1_89;
     wire data_out_1_89;

     reg pivot_in_1_89;
     wire pivot_out_1_89;

     always @(posedge clk) begin
         op_in_1_89 <= op_out_1_88;
         pivot_in_1_89 <= pivot_out_1_88;
         start_in_1_89 <= start_out_1_88;
     end

     always @(posedge clk) begin
         data_in_1_89 <= data_out_0_89;
     end
  
     processor_AB AB_1_89 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_89),
       .start_in   (start_in_1_89),
       .op_in      (op_in_1_89),
       .pivot_in   (pivot_in_1_89),
       .start_out  (start_out_1_89),
       .data_out   (data_out_1_89),
       .op_out     (op_out_1_89),
       .pivot_out  (pivot_out_1_89),
       .r          (r_1_89)
     );

  // row 1, col 90

     reg start_in_1_90;
     wire start_out_1_90;

     reg [1:0] op_in_1_90;
     wire [1:0] op_out_1_90;

     wire r_1_90;

     reg data_in_1_90;
     wire data_out_1_90;

     reg pivot_in_1_90;
     wire pivot_out_1_90;

     always @(posedge clk) begin
         op_in_1_90 <= op_out_1_89;
         pivot_in_1_90 <= pivot_out_1_89;
         start_in_1_90 <= start_out_1_89;
     end

     always @(posedge clk) begin
         data_in_1_90 <= data_out_0_90;
     end
  
     processor_AB AB_1_90 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_90),
       .start_in   (start_in_1_90),
       .op_in      (op_in_1_90),
       .pivot_in   (pivot_in_1_90),
       .start_out  (start_out_1_90),
       .data_out   (data_out_1_90),
       .op_out     (op_out_1_90),
       .pivot_out  (pivot_out_1_90),
       .r          (r_1_90)
     );

  // row 1, col 91

     reg start_in_1_91;
     wire start_out_1_91;

     reg [1:0] op_in_1_91;
     wire [1:0] op_out_1_91;

     wire r_1_91;

     reg data_in_1_91;
     wire data_out_1_91;

     reg pivot_in_1_91;
     wire pivot_out_1_91;

     always @(posedge clk) begin
         op_in_1_91 <= op_out_1_90;
         pivot_in_1_91 <= pivot_out_1_90;
         start_in_1_91 <= start_out_1_90;
     end

     always @(posedge clk) begin
         data_in_1_91 <= data_out_0_91;
     end
  
     processor_AB AB_1_91 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_91),
       .start_in   (start_in_1_91),
       .op_in      (op_in_1_91),
       .pivot_in   (pivot_in_1_91),
       .start_out  (start_out_1_91),
       .data_out   (data_out_1_91),
       .op_out     (op_out_1_91),
       .pivot_out  (pivot_out_1_91),
       .r          (r_1_91)
     );

  // row 1, col 92

     reg start_in_1_92;
     wire start_out_1_92;

     reg [1:0] op_in_1_92;
     wire [1:0] op_out_1_92;

     wire r_1_92;

     reg data_in_1_92;
     wire data_out_1_92;

     reg pivot_in_1_92;
     wire pivot_out_1_92;

     always @(posedge clk) begin
         op_in_1_92 <= op_out_1_91;
         pivot_in_1_92 <= pivot_out_1_91;
         start_in_1_92 <= start_out_1_91;
     end

     always @(posedge clk) begin
         data_in_1_92 <= data_out_0_92;
     end
  
     processor_AB AB_1_92 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_92),
       .start_in   (start_in_1_92),
       .op_in      (op_in_1_92),
       .pivot_in   (pivot_in_1_92),
       .start_out  (start_out_1_92),
       .data_out   (data_out_1_92),
       .op_out     (op_out_1_92),
       .pivot_out  (pivot_out_1_92),
       .r          (r_1_92)
     );

  // row 1, col 93

     reg start_in_1_93;
     wire start_out_1_93;

     reg [1:0] op_in_1_93;
     wire [1:0] op_out_1_93;

     wire r_1_93;

     reg data_in_1_93;
     wire data_out_1_93;

     reg pivot_in_1_93;
     wire pivot_out_1_93;

     always @(posedge clk) begin
         op_in_1_93 <= op_out_1_92;
         pivot_in_1_93 <= pivot_out_1_92;
         start_in_1_93 <= start_out_1_92;
     end

     always @(posedge clk) begin
         data_in_1_93 <= data_out_0_93;
     end
  
     processor_AB AB_1_93 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_93),
       .start_in   (start_in_1_93),
       .op_in      (op_in_1_93),
       .pivot_in   (pivot_in_1_93),
       .start_out  (start_out_1_93),
       .data_out   (data_out_1_93),
       .op_out     (op_out_1_93),
       .pivot_out  (pivot_out_1_93),
       .r          (r_1_93)
     );

  // row 1, col 94

     reg start_in_1_94;
     wire start_out_1_94;

     reg [1:0] op_in_1_94;
     wire [1:0] op_out_1_94;

     wire r_1_94;

     reg data_in_1_94;
     wire data_out_1_94;

     reg pivot_in_1_94;
     wire pivot_out_1_94;

     always @(posedge clk) begin
         op_in_1_94 <= op_out_1_93;
         pivot_in_1_94 <= pivot_out_1_93;
         start_in_1_94 <= start_out_1_93;
     end

     always @(posedge clk) begin
         data_in_1_94 <= data_out_0_94;
     end
  
     processor_AB AB_1_94 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_94),
       .start_in   (start_in_1_94),
       .op_in      (op_in_1_94),
       .pivot_in   (pivot_in_1_94),
       .start_out  (start_out_1_94),
       .data_out   (data_out_1_94),
       .op_out     (op_out_1_94),
       .pivot_out  (pivot_out_1_94),
       .r          (r_1_94)
     );

  // row 1, col 95

     reg start_in_1_95;
     wire start_out_1_95;

     reg [1:0] op_in_1_95;
     wire [1:0] op_out_1_95;

     wire r_1_95;

     reg data_in_1_95;
     wire data_out_1_95;

     reg pivot_in_1_95;
     wire pivot_out_1_95;

     always @(posedge clk) begin
         op_in_1_95 <= op_out_1_94;
         pivot_in_1_95 <= pivot_out_1_94;
         start_in_1_95 <= start_out_1_94;
     end

     always @(posedge clk) begin
         data_in_1_95 <= data_out_0_95;
     end
  
     processor_AB AB_1_95 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_95),
       .start_in   (start_in_1_95),
       .op_in      (op_in_1_95),
       .pivot_in   (pivot_in_1_95),
       .start_out  (start_out_1_95),
       .data_out   (data_out_1_95),
       .op_out     (op_out_1_95),
       .pivot_out  (pivot_out_1_95),
       .r          (r_1_95)
     );

  // row 1, col 96

     reg start_in_1_96;
     wire start_out_1_96;

     reg [1:0] op_in_1_96;
     wire [1:0] op_out_1_96;

     wire r_1_96;

     reg data_in_1_96;
     wire data_out_1_96;

     reg pivot_in_1_96;
     wire pivot_out_1_96;

     always @(posedge clk) begin
         op_in_1_96 <= op_out_1_95;
         pivot_in_1_96 <= pivot_out_1_95;
         start_in_1_96 <= start_out_1_95;
     end

     always @(posedge clk) begin
         data_in_1_96 <= data_out_0_96;
     end
  
     processor_AB AB_1_96 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_96),
       .start_in   (start_in_1_96),
       .op_in      (op_in_1_96),
       .pivot_in   (pivot_in_1_96),
       .start_out  (start_out_1_96),
       .data_out   (data_out_1_96),
       .op_out     (op_out_1_96),
       .pivot_out  (pivot_out_1_96),
       .r          (r_1_96)
     );

  // row 1, col 97

     reg start_in_1_97;
     wire start_out_1_97;

     reg [1:0] op_in_1_97;
     wire [1:0] op_out_1_97;

     wire r_1_97;

     reg data_in_1_97;
     wire data_out_1_97;

     reg pivot_in_1_97;
     wire pivot_out_1_97;

     always @(posedge clk) begin
         op_in_1_97 <= op_out_1_96;
         pivot_in_1_97 <= pivot_out_1_96;
         start_in_1_97 <= start_out_1_96;
     end

     always @(posedge clk) begin
         data_in_1_97 <= data_out_0_97;
     end
  
     processor_AB AB_1_97 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_97),
       .start_in   (start_in_1_97),
       .op_in      (op_in_1_97),
       .pivot_in   (pivot_in_1_97),
       .start_out  (start_out_1_97),
       .data_out   (data_out_1_97),
       .op_out     (op_out_1_97),
       .pivot_out  (pivot_out_1_97),
       .r          (r_1_97)
     );

  // row 1, col 98

     reg start_in_1_98;
     wire start_out_1_98;

     reg [1:0] op_in_1_98;
     wire [1:0] op_out_1_98;

     wire r_1_98;

     reg data_in_1_98;
     wire data_out_1_98;

     reg pivot_in_1_98;
     wire pivot_out_1_98;

     always @(posedge clk) begin
         op_in_1_98 <= op_out_1_97;
         pivot_in_1_98 <= pivot_out_1_97;
         start_in_1_98 <= start_out_1_97;
     end

     always @(posedge clk) begin
         data_in_1_98 <= data_out_0_98;
     end
  
     processor_AB AB_1_98 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_98),
       .start_in   (start_in_1_98),
       .op_in      (op_in_1_98),
       .pivot_in   (pivot_in_1_98),
       .start_out  (start_out_1_98),
       .data_out   (data_out_1_98),
       .op_out     (op_out_1_98),
       .pivot_out  (pivot_out_1_98),
       .r          (r_1_98)
     );

  // row 1, col 99

     reg start_in_1_99;
     wire start_out_1_99;

     reg [1:0] op_in_1_99;
     wire [1:0] op_out_1_99;

     wire r_1_99;

     reg data_in_1_99;
     wire data_out_1_99;

     reg pivot_in_1_99;
     wire pivot_out_1_99;

     always @(posedge clk) begin
         op_in_1_99 <= op_out_1_98;
         pivot_in_1_99 <= pivot_out_1_98;
         start_in_1_99 <= start_out_1_98;
     end

     always @(posedge clk) begin
         data_in_1_99 <= data_out_0_99;
     end
  
     processor_AB AB_1_99 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_99),
       .start_in   (start_in_1_99),
       .op_in      (op_in_1_99),
       .pivot_in   (pivot_in_1_99),
       .start_out  (start_out_1_99),
       .data_out   (data_out_1_99),
       .op_out     (op_out_1_99),
       .pivot_out  (pivot_out_1_99),
       .r          (r_1_99)
     );

  // row 1, col 100

     reg start_in_1_100;
     wire start_out_1_100;

     reg [1:0] op_in_1_100;
     wire [1:0] op_out_1_100;

     wire r_1_100;

     reg data_in_1_100;
     wire data_out_1_100;

     reg pivot_in_1_100;
     wire pivot_out_1_100;

     always @(posedge clk) begin
         op_in_1_100 <= op_out_1_99;
         pivot_in_1_100 <= pivot_out_1_99;
         start_in_1_100 <= start_out_1_99;
     end

     always @(posedge clk) begin
         data_in_1_100 <= data_out_0_100;
     end
  
     processor_AB AB_1_100 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_100),
       .start_in   (start_in_1_100),
       .op_in      (op_in_1_100),
       .pivot_in   (pivot_in_1_100),
       .start_out  (start_out_1_100),
       .data_out   (data_out_1_100),
       .op_out     (op_out_1_100),
       .pivot_out  (pivot_out_1_100),
       .r          (r_1_100)
     );

  /////////////////////////////////////
  // row 2
  // row 2, col 0

     wire start_in_2_0;
     wire start_out_2_0;

     wire [1:0] op_in_2_0;
     wire [1:0] op_out_2_0;

     wire r_2_0;

     reg data_in_2_0;
     wire data_out_2_0;

     wire pivot_in_2_0;
     wire pivout_out_2_0;

     assign op_in_2_0 = mode & start ? 2'b01 : 2'b00;
     assign pivot_in_2_0 = 0;

     assign start_in_2_0 = start_row[2]; 

     always @(posedge clk) begin
         data_in_2_0 <= data_out_1_0;
     end

     processor_AB AB_2_0 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_0),
       .start_in   (start_in_2_0),
       .op_in      (op_in_2_0),
       .pivot_in   (pivot_in_2_0),
       .start_out  (start_out_2_0),
       .data_out   (data_out_2_0),
       .op_out     (op_out_2_0),
       .pivot_out  (pivot_out_2_0),
       .r          (r_2_0)
     );

  // row 2, col 1

     reg start_in_2_1;
     wire start_out_2_1;

     reg [1:0] op_in_2_1;
     wire [1:0] op_out_2_1;

     wire r_2_1;

     reg data_in_2_1;
     wire data_out_2_1;

     reg pivot_in_2_1;
     wire pivot_out_2_1;

     always @(posedge clk) begin
         op_in_2_1 <= op_out_2_0;
         pivot_in_2_1 <= pivot_out_2_0;
         start_in_2_1 <= start_out_2_0;
     end

     always @(posedge clk) begin
         data_in_2_1 <= data_out_1_1;
     end
  
     processor_AB AB_2_1 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_1),
       .start_in   (start_in_2_1),
       .op_in      (op_in_2_1),
       .pivot_in   (pivot_in_2_1),
       .start_out  (start_out_2_1),
       .data_out   (data_out_2_1),
       .op_out     (op_out_2_1),
       .pivot_out  (pivot_out_2_1),
       .r          (r_2_1)
     );

  // row 2, col 2

     reg start_in_2_2;
     wire start_out_2_2;

     reg [1:0] op_in_2_2;
     wire [1:0] op_out_2_2;

     wire r_2_2;

     reg data_in_2_2;
     wire data_out_2_2;

     reg pivot_in_2_2;
     wire pivot_out_2_2;

     always @(posedge clk) begin
         op_in_2_2 <= op_out_2_1;
         pivot_in_2_2 <= pivot_out_2_1;
         start_in_2_2 <= start_out_2_1;
     end

     always @(posedge clk) begin
         data_in_2_2 <= data_out_1_2;
     end
  
     processor_AB AB_2_2 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_2),
       .start_in   (start_in_2_2),
       .op_in      (op_in_2_2),
       .pivot_in   (pivot_in_2_2),
       .start_out  (start_out_2_2),
       .data_out   (data_out_2_2),
       .op_out     (op_out_2_2),
       .pivot_out  (pivot_out_2_2),
       .r          (r_2_2)
     );

  // row 2, col 3

     reg start_in_2_3;
     wire start_out_2_3;

     reg [1:0] op_in_2_3;
     wire [1:0] op_out_2_3;

     wire r_2_3;

     reg data_in_2_3;
     wire data_out_2_3;

     reg pivot_in_2_3;
     wire pivot_out_2_3;

     always @(posedge clk) begin
         op_in_2_3 <= op_out_2_2;
         pivot_in_2_3 <= pivot_out_2_2;
         start_in_2_3 <= start_out_2_2;
     end

     always @(posedge clk) begin
         data_in_2_3 <= data_out_1_3;
     end
  
     processor_AB AB_2_3 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_3),
       .start_in   (start_in_2_3),
       .op_in      (op_in_2_3),
       .pivot_in   (pivot_in_2_3),
       .start_out  (start_out_2_3),
       .data_out   (data_out_2_3),
       .op_out     (op_out_2_3),
       .pivot_out  (pivot_out_2_3),
       .r          (r_2_3)
     );

  // row 2, col 4

     reg start_in_2_4;
     wire start_out_2_4;

     reg [1:0] op_in_2_4;
     wire [1:0] op_out_2_4;

     wire r_2_4;

     reg data_in_2_4;
     wire data_out_2_4;

     reg pivot_in_2_4;
     wire pivot_out_2_4;

     always @(posedge clk) begin
         op_in_2_4 <= op_out_2_3;
         pivot_in_2_4 <= pivot_out_2_3;
         start_in_2_4 <= start_out_2_3;
     end

     always @(posedge clk) begin
         data_in_2_4 <= data_out_1_4;
     end
  
     processor_AB AB_2_4 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_4),
       .start_in   (start_in_2_4),
       .op_in      (op_in_2_4),
       .pivot_in   (pivot_in_2_4),
       .start_out  (start_out_2_4),
       .data_out   (data_out_2_4),
       .op_out     (op_out_2_4),
       .pivot_out  (pivot_out_2_4),
       .r          (r_2_4)
     );

  // row 2, col 5

     reg start_in_2_5;
     wire start_out_2_5;

     reg [1:0] op_in_2_5;
     wire [1:0] op_out_2_5;

     wire r_2_5;

     reg data_in_2_5;
     wire data_out_2_5;

     reg pivot_in_2_5;
     wire pivot_out_2_5;

     always @(posedge clk) begin
         op_in_2_5 <= op_out_2_4;
         pivot_in_2_5 <= pivot_out_2_4;
         start_in_2_5 <= start_out_2_4;
     end

     always @(posedge clk) begin
         data_in_2_5 <= data_out_1_5;
     end
  
     processor_AB AB_2_5 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_5),
       .start_in   (start_in_2_5),
       .op_in      (op_in_2_5),
       .pivot_in   (pivot_in_2_5),
       .start_out  (start_out_2_5),
       .data_out   (data_out_2_5),
       .op_out     (op_out_2_5),
       .pivot_out  (pivot_out_2_5),
       .r          (r_2_5)
     );

  // row 2, col 6

     reg start_in_2_6;
     wire start_out_2_6;

     reg [1:0] op_in_2_6;
     wire [1:0] op_out_2_6;

     wire r_2_6;

     reg data_in_2_6;
     wire data_out_2_6;

     reg pivot_in_2_6;
     wire pivot_out_2_6;

     always @(posedge clk) begin
         op_in_2_6 <= op_out_2_5;
         pivot_in_2_6 <= pivot_out_2_5;
         start_in_2_6 <= start_out_2_5;
     end

     always @(posedge clk) begin
         data_in_2_6 <= data_out_1_6;
     end
  
     processor_AB AB_2_6 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_6),
       .start_in   (start_in_2_6),
       .op_in      (op_in_2_6),
       .pivot_in   (pivot_in_2_6),
       .start_out  (start_out_2_6),
       .data_out   (data_out_2_6),
       .op_out     (op_out_2_6),
       .pivot_out  (pivot_out_2_6),
       .r          (r_2_6)
     );

  // row 2, col 7

     reg start_in_2_7;
     wire start_out_2_7;

     reg [1:0] op_in_2_7;
     wire [1:0] op_out_2_7;

     wire r_2_7;

     reg data_in_2_7;
     wire data_out_2_7;

     reg pivot_in_2_7;
     wire pivot_out_2_7;

     always @(posedge clk) begin
         op_in_2_7 <= op_out_2_6;
         pivot_in_2_7 <= pivot_out_2_6;
         start_in_2_7 <= start_out_2_6;
     end

     always @(posedge clk) begin
         data_in_2_7 <= data_out_1_7;
     end
  
     processor_AB AB_2_7 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_7),
       .start_in   (start_in_2_7),
       .op_in      (op_in_2_7),
       .pivot_in   (pivot_in_2_7),
       .start_out  (start_out_2_7),
       .data_out   (data_out_2_7),
       .op_out     (op_out_2_7),
       .pivot_out  (pivot_out_2_7),
       .r          (r_2_7)
     );

  // row 2, col 8

     reg start_in_2_8;
     wire start_out_2_8;

     reg [1:0] op_in_2_8;
     wire [1:0] op_out_2_8;

     wire r_2_8;

     reg data_in_2_8;
     wire data_out_2_8;

     reg pivot_in_2_8;
     wire pivot_out_2_8;

     always @(posedge clk) begin
         op_in_2_8 <= op_out_2_7;
         pivot_in_2_8 <= pivot_out_2_7;
         start_in_2_8 <= start_out_2_7;
     end

     always @(posedge clk) begin
         data_in_2_8 <= data_out_1_8;
     end
  
     processor_AB AB_2_8 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_8),
       .start_in   (start_in_2_8),
       .op_in      (op_in_2_8),
       .pivot_in   (pivot_in_2_8),
       .start_out  (start_out_2_8),
       .data_out   (data_out_2_8),
       .op_out     (op_out_2_8),
       .pivot_out  (pivot_out_2_8),
       .r          (r_2_8)
     );

  // row 2, col 9

     reg start_in_2_9;
     wire start_out_2_9;

     reg [1:0] op_in_2_9;
     wire [1:0] op_out_2_9;

     wire r_2_9;

     reg data_in_2_9;
     wire data_out_2_9;

     reg pivot_in_2_9;
     wire pivot_out_2_9;

     always @(posedge clk) begin
         op_in_2_9 <= op_out_2_8;
         pivot_in_2_9 <= pivot_out_2_8;
         start_in_2_9 <= start_out_2_8;
     end

     always @(posedge clk) begin
         data_in_2_9 <= data_out_1_9;
     end
  
     processor_AB AB_2_9 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_9),
       .start_in   (start_in_2_9),
       .op_in      (op_in_2_9),
       .pivot_in   (pivot_in_2_9),
       .start_out  (start_out_2_9),
       .data_out   (data_out_2_9),
       .op_out     (op_out_2_9),
       .pivot_out  (pivot_out_2_9),
       .r          (r_2_9)
     );

  // row 2, col 10

     reg start_in_2_10;
     wire start_out_2_10;

     reg [1:0] op_in_2_10;
     wire [1:0] op_out_2_10;

     wire r_2_10;

     reg data_in_2_10;
     wire data_out_2_10;

     reg pivot_in_2_10;
     wire pivot_out_2_10;

     always @(posedge clk) begin
         op_in_2_10 <= op_out_2_9;
         pivot_in_2_10 <= pivot_out_2_9;
         start_in_2_10 <= start_out_2_9;
     end

     always @(posedge clk) begin
         data_in_2_10 <= data_out_1_10;
     end
  
     processor_AB AB_2_10 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_10),
       .start_in   (start_in_2_10),
       .op_in      (op_in_2_10),
       .pivot_in   (pivot_in_2_10),
       .start_out  (start_out_2_10),
       .data_out   (data_out_2_10),
       .op_out     (op_out_2_10),
       .pivot_out  (pivot_out_2_10),
       .r          (r_2_10)
     );

  // row 2, col 11

     reg start_in_2_11;
     wire start_out_2_11;

     reg [1:0] op_in_2_11;
     wire [1:0] op_out_2_11;

     wire r_2_11;

     reg data_in_2_11;
     wire data_out_2_11;

     reg pivot_in_2_11;
     wire pivot_out_2_11;

     always @(posedge clk) begin
         op_in_2_11 <= op_out_2_10;
         pivot_in_2_11 <= pivot_out_2_10;
         start_in_2_11 <= start_out_2_10;
     end

     always @(posedge clk) begin
         data_in_2_11 <= data_out_1_11;
     end
  
     processor_AB AB_2_11 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_11),
       .start_in   (start_in_2_11),
       .op_in      (op_in_2_11),
       .pivot_in   (pivot_in_2_11),
       .start_out  (start_out_2_11),
       .data_out   (data_out_2_11),
       .op_out     (op_out_2_11),
       .pivot_out  (pivot_out_2_11),
       .r          (r_2_11)
     );

  // row 2, col 12

     reg start_in_2_12;
     wire start_out_2_12;

     reg [1:0] op_in_2_12;
     wire [1:0] op_out_2_12;

     wire r_2_12;

     reg data_in_2_12;
     wire data_out_2_12;

     reg pivot_in_2_12;
     wire pivot_out_2_12;

     always @(posedge clk) begin
         op_in_2_12 <= op_out_2_11;
         pivot_in_2_12 <= pivot_out_2_11;
         start_in_2_12 <= start_out_2_11;
     end

     always @(posedge clk) begin
         data_in_2_12 <= data_out_1_12;
     end
  
     processor_AB AB_2_12 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_12),
       .start_in   (start_in_2_12),
       .op_in      (op_in_2_12),
       .pivot_in   (pivot_in_2_12),
       .start_out  (start_out_2_12),
       .data_out   (data_out_2_12),
       .op_out     (op_out_2_12),
       .pivot_out  (pivot_out_2_12),
       .r          (r_2_12)
     );

  // row 2, col 13

     reg start_in_2_13;
     wire start_out_2_13;

     reg [1:0] op_in_2_13;
     wire [1:0] op_out_2_13;

     wire r_2_13;

     reg data_in_2_13;
     wire data_out_2_13;

     reg pivot_in_2_13;
     wire pivot_out_2_13;

     always @(posedge clk) begin
         op_in_2_13 <= op_out_2_12;
         pivot_in_2_13 <= pivot_out_2_12;
         start_in_2_13 <= start_out_2_12;
     end

     always @(posedge clk) begin
         data_in_2_13 <= data_out_1_13;
     end
  
     processor_AB AB_2_13 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_13),
       .start_in   (start_in_2_13),
       .op_in      (op_in_2_13),
       .pivot_in   (pivot_in_2_13),
       .start_out  (start_out_2_13),
       .data_out   (data_out_2_13),
       .op_out     (op_out_2_13),
       .pivot_out  (pivot_out_2_13),
       .r          (r_2_13)
     );

  // row 2, col 14

     reg start_in_2_14;
     wire start_out_2_14;

     reg [1:0] op_in_2_14;
     wire [1:0] op_out_2_14;

     wire r_2_14;

     reg data_in_2_14;
     wire data_out_2_14;

     reg pivot_in_2_14;
     wire pivot_out_2_14;

     always @(posedge clk) begin
         op_in_2_14 <= op_out_2_13;
         pivot_in_2_14 <= pivot_out_2_13;
         start_in_2_14 <= start_out_2_13;
     end

     always @(posedge clk) begin
         data_in_2_14 <= data_out_1_14;
     end
  
     processor_AB AB_2_14 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_14),
       .start_in   (start_in_2_14),
       .op_in      (op_in_2_14),
       .pivot_in   (pivot_in_2_14),
       .start_out  (start_out_2_14),
       .data_out   (data_out_2_14),
       .op_out     (op_out_2_14),
       .pivot_out  (pivot_out_2_14),
       .r          (r_2_14)
     );

  // row 2, col 15

     reg start_in_2_15;
     wire start_out_2_15;

     reg [1:0] op_in_2_15;
     wire [1:0] op_out_2_15;

     wire r_2_15;

     reg data_in_2_15;
     wire data_out_2_15;

     reg pivot_in_2_15;
     wire pivot_out_2_15;

     always @(posedge clk) begin
         op_in_2_15 <= op_out_2_14;
         pivot_in_2_15 <= pivot_out_2_14;
         start_in_2_15 <= start_out_2_14;
     end

     always @(posedge clk) begin
         data_in_2_15 <= data_out_1_15;
     end
  
     processor_AB AB_2_15 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_15),
       .start_in   (start_in_2_15),
       .op_in      (op_in_2_15),
       .pivot_in   (pivot_in_2_15),
       .start_out  (start_out_2_15),
       .data_out   (data_out_2_15),
       .op_out     (op_out_2_15),
       .pivot_out  (pivot_out_2_15),
       .r          (r_2_15)
     );

  // row 2, col 16

     reg start_in_2_16;
     wire start_out_2_16;

     reg [1:0] op_in_2_16;
     wire [1:0] op_out_2_16;

     wire r_2_16;

     reg data_in_2_16;
     wire data_out_2_16;

     reg pivot_in_2_16;
     wire pivot_out_2_16;

     always @(posedge clk) begin
         op_in_2_16 <= op_out_2_15;
         pivot_in_2_16 <= pivot_out_2_15;
         start_in_2_16 <= start_out_2_15;
     end

     always @(posedge clk) begin
         data_in_2_16 <= data_out_1_16;
     end
  
     processor_AB AB_2_16 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_16),
       .start_in   (start_in_2_16),
       .op_in      (op_in_2_16),
       .pivot_in   (pivot_in_2_16),
       .start_out  (start_out_2_16),
       .data_out   (data_out_2_16),
       .op_out     (op_out_2_16),
       .pivot_out  (pivot_out_2_16),
       .r          (r_2_16)
     );

  // row 2, col 17

     reg start_in_2_17;
     wire start_out_2_17;

     reg [1:0] op_in_2_17;
     wire [1:0] op_out_2_17;

     wire r_2_17;

     reg data_in_2_17;
     wire data_out_2_17;

     reg pivot_in_2_17;
     wire pivot_out_2_17;

     always @(posedge clk) begin
         op_in_2_17 <= op_out_2_16;
         pivot_in_2_17 <= pivot_out_2_16;
         start_in_2_17 <= start_out_2_16;
     end

     always @(posedge clk) begin
         data_in_2_17 <= data_out_1_17;
     end
  
     processor_AB AB_2_17 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_17),
       .start_in   (start_in_2_17),
       .op_in      (op_in_2_17),
       .pivot_in   (pivot_in_2_17),
       .start_out  (start_out_2_17),
       .data_out   (data_out_2_17),
       .op_out     (op_out_2_17),
       .pivot_out  (pivot_out_2_17),
       .r          (r_2_17)
     );

  // row 2, col 18

     reg start_in_2_18;
     wire start_out_2_18;

     reg [1:0] op_in_2_18;
     wire [1:0] op_out_2_18;

     wire r_2_18;

     reg data_in_2_18;
     wire data_out_2_18;

     reg pivot_in_2_18;
     wire pivot_out_2_18;

     always @(posedge clk) begin
         op_in_2_18 <= op_out_2_17;
         pivot_in_2_18 <= pivot_out_2_17;
         start_in_2_18 <= start_out_2_17;
     end

     always @(posedge clk) begin
         data_in_2_18 <= data_out_1_18;
     end
  
     processor_AB AB_2_18 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_18),
       .start_in   (start_in_2_18),
       .op_in      (op_in_2_18),
       .pivot_in   (pivot_in_2_18),
       .start_out  (start_out_2_18),
       .data_out   (data_out_2_18),
       .op_out     (op_out_2_18),
       .pivot_out  (pivot_out_2_18),
       .r          (r_2_18)
     );

  // row 2, col 19

     reg start_in_2_19;
     wire start_out_2_19;

     reg [1:0] op_in_2_19;
     wire [1:0] op_out_2_19;

     wire r_2_19;

     reg data_in_2_19;
     wire data_out_2_19;

     reg pivot_in_2_19;
     wire pivot_out_2_19;

     always @(posedge clk) begin
         op_in_2_19 <= op_out_2_18;
         pivot_in_2_19 <= pivot_out_2_18;
         start_in_2_19 <= start_out_2_18;
     end

     always @(posedge clk) begin
         data_in_2_19 <= data_out_1_19;
     end
  
     processor_AB AB_2_19 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_19),
       .start_in   (start_in_2_19),
       .op_in      (op_in_2_19),
       .pivot_in   (pivot_in_2_19),
       .start_out  (start_out_2_19),
       .data_out   (data_out_2_19),
       .op_out     (op_out_2_19),
       .pivot_out  (pivot_out_2_19),
       .r          (r_2_19)
     );

  // row 2, col 20

     reg start_in_2_20;
     wire start_out_2_20;

     reg [1:0] op_in_2_20;
     wire [1:0] op_out_2_20;

     wire r_2_20;

     reg data_in_2_20;
     wire data_out_2_20;

     reg pivot_in_2_20;
     wire pivot_out_2_20;

     always @(posedge clk) begin
         op_in_2_20 <= op_out_2_19;
         pivot_in_2_20 <= pivot_out_2_19;
         start_in_2_20 <= start_out_2_19;
     end

     always @(posedge clk) begin
         data_in_2_20 <= data_out_1_20;
     end
  
     processor_AB AB_2_20 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_20),
       .start_in   (start_in_2_20),
       .op_in      (op_in_2_20),
       .pivot_in   (pivot_in_2_20),
       .start_out  (start_out_2_20),
       .data_out   (data_out_2_20),
       .op_out     (op_out_2_20),
       .pivot_out  (pivot_out_2_20),
       .r          (r_2_20)
     );

  // row 2, col 21

     reg start_in_2_21;
     wire start_out_2_21;

     reg [1:0] op_in_2_21;
     wire [1:0] op_out_2_21;

     wire r_2_21;

     reg data_in_2_21;
     wire data_out_2_21;

     reg pivot_in_2_21;
     wire pivot_out_2_21;

     always @(posedge clk) begin
         op_in_2_21 <= op_out_2_20;
         pivot_in_2_21 <= pivot_out_2_20;
         start_in_2_21 <= start_out_2_20;
     end

     always @(posedge clk) begin
         data_in_2_21 <= data_out_1_21;
     end
  
     processor_AB AB_2_21 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_21),
       .start_in   (start_in_2_21),
       .op_in      (op_in_2_21),
       .pivot_in   (pivot_in_2_21),
       .start_out  (start_out_2_21),
       .data_out   (data_out_2_21),
       .op_out     (op_out_2_21),
       .pivot_out  (pivot_out_2_21),
       .r          (r_2_21)
     );

  // row 2, col 22

     reg start_in_2_22;
     wire start_out_2_22;

     reg [1:0] op_in_2_22;
     wire [1:0] op_out_2_22;

     wire r_2_22;

     reg data_in_2_22;
     wire data_out_2_22;

     reg pivot_in_2_22;
     wire pivot_out_2_22;

     always @(posedge clk) begin
         op_in_2_22 <= op_out_2_21;
         pivot_in_2_22 <= pivot_out_2_21;
         start_in_2_22 <= start_out_2_21;
     end

     always @(posedge clk) begin
         data_in_2_22 <= data_out_1_22;
     end
  
     processor_AB AB_2_22 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_22),
       .start_in   (start_in_2_22),
       .op_in      (op_in_2_22),
       .pivot_in   (pivot_in_2_22),
       .start_out  (start_out_2_22),
       .data_out   (data_out_2_22),
       .op_out     (op_out_2_22),
       .pivot_out  (pivot_out_2_22),
       .r          (r_2_22)
     );

  // row 2, col 23

     reg start_in_2_23;
     wire start_out_2_23;

     reg [1:0] op_in_2_23;
     wire [1:0] op_out_2_23;

     wire r_2_23;

     reg data_in_2_23;
     wire data_out_2_23;

     reg pivot_in_2_23;
     wire pivot_out_2_23;

     always @(posedge clk) begin
         op_in_2_23 <= op_out_2_22;
         pivot_in_2_23 <= pivot_out_2_22;
         start_in_2_23 <= start_out_2_22;
     end

     always @(posedge clk) begin
         data_in_2_23 <= data_out_1_23;
     end
  
     processor_AB AB_2_23 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_23),
       .start_in   (start_in_2_23),
       .op_in      (op_in_2_23),
       .pivot_in   (pivot_in_2_23),
       .start_out  (start_out_2_23),
       .data_out   (data_out_2_23),
       .op_out     (op_out_2_23),
       .pivot_out  (pivot_out_2_23),
       .r          (r_2_23)
     );

  // row 2, col 24

     reg start_in_2_24;
     wire start_out_2_24;

     reg [1:0] op_in_2_24;
     wire [1:0] op_out_2_24;

     wire r_2_24;

     reg data_in_2_24;
     wire data_out_2_24;

     reg pivot_in_2_24;
     wire pivot_out_2_24;

     always @(posedge clk) begin
         op_in_2_24 <= op_out_2_23;
         pivot_in_2_24 <= pivot_out_2_23;
         start_in_2_24 <= start_out_2_23;
     end

     always @(posedge clk) begin
         data_in_2_24 <= data_out_1_24;
     end
  
     processor_AB AB_2_24 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_24),
       .start_in   (start_in_2_24),
       .op_in      (op_in_2_24),
       .pivot_in   (pivot_in_2_24),
       .start_out  (start_out_2_24),
       .data_out   (data_out_2_24),
       .op_out     (op_out_2_24),
       .pivot_out  (pivot_out_2_24),
       .r          (r_2_24)
     );

  // row 2, col 25

     reg start_in_2_25;
     wire start_out_2_25;

     reg [1:0] op_in_2_25;
     wire [1:0] op_out_2_25;

     wire r_2_25;

     reg data_in_2_25;
     wire data_out_2_25;

     reg pivot_in_2_25;
     wire pivot_out_2_25;

     always @(posedge clk) begin
         op_in_2_25 <= op_out_2_24;
         pivot_in_2_25 <= pivot_out_2_24;
         start_in_2_25 <= start_out_2_24;
     end

     always @(posedge clk) begin
         data_in_2_25 <= data_out_1_25;
     end
  
     processor_AB AB_2_25 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_25),
       .start_in   (start_in_2_25),
       .op_in      (op_in_2_25),
       .pivot_in   (pivot_in_2_25),
       .start_out  (start_out_2_25),
       .data_out   (data_out_2_25),
       .op_out     (op_out_2_25),
       .pivot_out  (pivot_out_2_25),
       .r          (r_2_25)
     );

  // row 2, col 26

     reg start_in_2_26;
     wire start_out_2_26;

     reg [1:0] op_in_2_26;
     wire [1:0] op_out_2_26;

     wire r_2_26;

     reg data_in_2_26;
     wire data_out_2_26;

     reg pivot_in_2_26;
     wire pivot_out_2_26;

     always @(posedge clk) begin
         op_in_2_26 <= op_out_2_25;
         pivot_in_2_26 <= pivot_out_2_25;
         start_in_2_26 <= start_out_2_25;
     end

     always @(posedge clk) begin
         data_in_2_26 <= data_out_1_26;
     end
  
     processor_AB AB_2_26 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_26),
       .start_in   (start_in_2_26),
       .op_in      (op_in_2_26),
       .pivot_in   (pivot_in_2_26),
       .start_out  (start_out_2_26),
       .data_out   (data_out_2_26),
       .op_out     (op_out_2_26),
       .pivot_out  (pivot_out_2_26),
       .r          (r_2_26)
     );

  // row 2, col 27

     reg start_in_2_27;
     wire start_out_2_27;

     reg [1:0] op_in_2_27;
     wire [1:0] op_out_2_27;

     wire r_2_27;

     reg data_in_2_27;
     wire data_out_2_27;

     reg pivot_in_2_27;
     wire pivot_out_2_27;

     always @(posedge clk) begin
         op_in_2_27 <= op_out_2_26;
         pivot_in_2_27 <= pivot_out_2_26;
         start_in_2_27 <= start_out_2_26;
     end

     always @(posedge clk) begin
         data_in_2_27 <= data_out_1_27;
     end
  
     processor_AB AB_2_27 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_27),
       .start_in   (start_in_2_27),
       .op_in      (op_in_2_27),
       .pivot_in   (pivot_in_2_27),
       .start_out  (start_out_2_27),
       .data_out   (data_out_2_27),
       .op_out     (op_out_2_27),
       .pivot_out  (pivot_out_2_27),
       .r          (r_2_27)
     );

  // row 2, col 28

     reg start_in_2_28;
     wire start_out_2_28;

     reg [1:0] op_in_2_28;
     wire [1:0] op_out_2_28;

     wire r_2_28;

     reg data_in_2_28;
     wire data_out_2_28;

     reg pivot_in_2_28;
     wire pivot_out_2_28;

     always @(posedge clk) begin
         op_in_2_28 <= op_out_2_27;
         pivot_in_2_28 <= pivot_out_2_27;
         start_in_2_28 <= start_out_2_27;
     end

     always @(posedge clk) begin
         data_in_2_28 <= data_out_1_28;
     end
  
     processor_AB AB_2_28 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_28),
       .start_in   (start_in_2_28),
       .op_in      (op_in_2_28),
       .pivot_in   (pivot_in_2_28),
       .start_out  (start_out_2_28),
       .data_out   (data_out_2_28),
       .op_out     (op_out_2_28),
       .pivot_out  (pivot_out_2_28),
       .r          (r_2_28)
     );

  // row 2, col 29

     reg start_in_2_29;
     wire start_out_2_29;

     reg [1:0] op_in_2_29;
     wire [1:0] op_out_2_29;

     wire r_2_29;

     reg data_in_2_29;
     wire data_out_2_29;

     reg pivot_in_2_29;
     wire pivot_out_2_29;

     always @(posedge clk) begin
         op_in_2_29 <= op_out_2_28;
         pivot_in_2_29 <= pivot_out_2_28;
         start_in_2_29 <= start_out_2_28;
     end

     always @(posedge clk) begin
         data_in_2_29 <= data_out_1_29;
     end
  
     processor_AB AB_2_29 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_29),
       .start_in   (start_in_2_29),
       .op_in      (op_in_2_29),
       .pivot_in   (pivot_in_2_29),
       .start_out  (start_out_2_29),
       .data_out   (data_out_2_29),
       .op_out     (op_out_2_29),
       .pivot_out  (pivot_out_2_29),
       .r          (r_2_29)
     );

  // row 2, col 30

     reg start_in_2_30;
     wire start_out_2_30;

     reg [1:0] op_in_2_30;
     wire [1:0] op_out_2_30;

     wire r_2_30;

     reg data_in_2_30;
     wire data_out_2_30;

     reg pivot_in_2_30;
     wire pivot_out_2_30;

     always @(posedge clk) begin
         op_in_2_30 <= op_out_2_29;
         pivot_in_2_30 <= pivot_out_2_29;
         start_in_2_30 <= start_out_2_29;
     end

     always @(posedge clk) begin
         data_in_2_30 <= data_out_1_30;
     end
  
     processor_AB AB_2_30 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_30),
       .start_in   (start_in_2_30),
       .op_in      (op_in_2_30),
       .pivot_in   (pivot_in_2_30),
       .start_out  (start_out_2_30),
       .data_out   (data_out_2_30),
       .op_out     (op_out_2_30),
       .pivot_out  (pivot_out_2_30),
       .r          (r_2_30)
     );

  // row 2, col 31

     reg start_in_2_31;
     wire start_out_2_31;

     reg [1:0] op_in_2_31;
     wire [1:0] op_out_2_31;

     wire r_2_31;

     reg data_in_2_31;
     wire data_out_2_31;

     reg pivot_in_2_31;
     wire pivot_out_2_31;

     always @(posedge clk) begin
         op_in_2_31 <= op_out_2_30;
         pivot_in_2_31 <= pivot_out_2_30;
         start_in_2_31 <= start_out_2_30;
     end

     always @(posedge clk) begin
         data_in_2_31 <= data_out_1_31;
     end
  
     processor_AB AB_2_31 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_31),
       .start_in   (start_in_2_31),
       .op_in      (op_in_2_31),
       .pivot_in   (pivot_in_2_31),
       .start_out  (start_out_2_31),
       .data_out   (data_out_2_31),
       .op_out     (op_out_2_31),
       .pivot_out  (pivot_out_2_31),
       .r          (r_2_31)
     );

  // row 2, col 32

     reg start_in_2_32;
     wire start_out_2_32;

     reg [1:0] op_in_2_32;
     wire [1:0] op_out_2_32;

     wire r_2_32;

     reg data_in_2_32;
     wire data_out_2_32;

     reg pivot_in_2_32;
     wire pivot_out_2_32;

     always @(posedge clk) begin
         op_in_2_32 <= op_out_2_31;
         pivot_in_2_32 <= pivot_out_2_31;
         start_in_2_32 <= start_out_2_31;
     end

     always @(posedge clk) begin
         data_in_2_32 <= data_out_1_32;
     end
  
     processor_AB AB_2_32 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_32),
       .start_in   (start_in_2_32),
       .op_in      (op_in_2_32),
       .pivot_in   (pivot_in_2_32),
       .start_out  (start_out_2_32),
       .data_out   (data_out_2_32),
       .op_out     (op_out_2_32),
       .pivot_out  (pivot_out_2_32),
       .r          (r_2_32)
     );

  // row 2, col 33

     reg start_in_2_33;
     wire start_out_2_33;

     reg [1:0] op_in_2_33;
     wire [1:0] op_out_2_33;

     wire r_2_33;

     reg data_in_2_33;
     wire data_out_2_33;

     reg pivot_in_2_33;
     wire pivot_out_2_33;

     always @(posedge clk) begin
         op_in_2_33 <= op_out_2_32;
         pivot_in_2_33 <= pivot_out_2_32;
         start_in_2_33 <= start_out_2_32;
     end

     always @(posedge clk) begin
         data_in_2_33 <= data_out_1_33;
     end
  
     processor_AB AB_2_33 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_33),
       .start_in   (start_in_2_33),
       .op_in      (op_in_2_33),
       .pivot_in   (pivot_in_2_33),
       .start_out  (start_out_2_33),
       .data_out   (data_out_2_33),
       .op_out     (op_out_2_33),
       .pivot_out  (pivot_out_2_33),
       .r          (r_2_33)
     );

  // row 2, col 34

     reg start_in_2_34;
     wire start_out_2_34;

     reg [1:0] op_in_2_34;
     wire [1:0] op_out_2_34;

     wire r_2_34;

     reg data_in_2_34;
     wire data_out_2_34;

     reg pivot_in_2_34;
     wire pivot_out_2_34;

     always @(posedge clk) begin
         op_in_2_34 <= op_out_2_33;
         pivot_in_2_34 <= pivot_out_2_33;
         start_in_2_34 <= start_out_2_33;
     end

     always @(posedge clk) begin
         data_in_2_34 <= data_out_1_34;
     end
  
     processor_AB AB_2_34 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_34),
       .start_in   (start_in_2_34),
       .op_in      (op_in_2_34),
       .pivot_in   (pivot_in_2_34),
       .start_out  (start_out_2_34),
       .data_out   (data_out_2_34),
       .op_out     (op_out_2_34),
       .pivot_out  (pivot_out_2_34),
       .r          (r_2_34)
     );

  // row 2, col 35

     reg start_in_2_35;
     wire start_out_2_35;

     reg [1:0] op_in_2_35;
     wire [1:0] op_out_2_35;

     wire r_2_35;

     reg data_in_2_35;
     wire data_out_2_35;

     reg pivot_in_2_35;
     wire pivot_out_2_35;

     always @(posedge clk) begin
         op_in_2_35 <= op_out_2_34;
         pivot_in_2_35 <= pivot_out_2_34;
         start_in_2_35 <= start_out_2_34;
     end

     always @(posedge clk) begin
         data_in_2_35 <= data_out_1_35;
     end
  
     processor_AB AB_2_35 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_35),
       .start_in   (start_in_2_35),
       .op_in      (op_in_2_35),
       .pivot_in   (pivot_in_2_35),
       .start_out  (start_out_2_35),
       .data_out   (data_out_2_35),
       .op_out     (op_out_2_35),
       .pivot_out  (pivot_out_2_35),
       .r          (r_2_35)
     );

  // row 2, col 36

     reg start_in_2_36;
     wire start_out_2_36;

     reg [1:0] op_in_2_36;
     wire [1:0] op_out_2_36;

     wire r_2_36;

     reg data_in_2_36;
     wire data_out_2_36;

     reg pivot_in_2_36;
     wire pivot_out_2_36;

     always @(posedge clk) begin
         op_in_2_36 <= op_out_2_35;
         pivot_in_2_36 <= pivot_out_2_35;
         start_in_2_36 <= start_out_2_35;
     end

     always @(posedge clk) begin
         data_in_2_36 <= data_out_1_36;
     end
  
     processor_AB AB_2_36 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_36),
       .start_in   (start_in_2_36),
       .op_in      (op_in_2_36),
       .pivot_in   (pivot_in_2_36),
       .start_out  (start_out_2_36),
       .data_out   (data_out_2_36),
       .op_out     (op_out_2_36),
       .pivot_out  (pivot_out_2_36),
       .r          (r_2_36)
     );

  // row 2, col 37

     reg start_in_2_37;
     wire start_out_2_37;

     reg [1:0] op_in_2_37;
     wire [1:0] op_out_2_37;

     wire r_2_37;

     reg data_in_2_37;
     wire data_out_2_37;

     reg pivot_in_2_37;
     wire pivot_out_2_37;

     always @(posedge clk) begin
         op_in_2_37 <= op_out_2_36;
         pivot_in_2_37 <= pivot_out_2_36;
         start_in_2_37 <= start_out_2_36;
     end

     always @(posedge clk) begin
         data_in_2_37 <= data_out_1_37;
     end
  
     processor_AB AB_2_37 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_37),
       .start_in   (start_in_2_37),
       .op_in      (op_in_2_37),
       .pivot_in   (pivot_in_2_37),
       .start_out  (start_out_2_37),
       .data_out   (data_out_2_37),
       .op_out     (op_out_2_37),
       .pivot_out  (pivot_out_2_37),
       .r          (r_2_37)
     );

  // row 2, col 38

     reg start_in_2_38;
     wire start_out_2_38;

     reg [1:0] op_in_2_38;
     wire [1:0] op_out_2_38;

     wire r_2_38;

     reg data_in_2_38;
     wire data_out_2_38;

     reg pivot_in_2_38;
     wire pivot_out_2_38;

     always @(posedge clk) begin
         op_in_2_38 <= op_out_2_37;
         pivot_in_2_38 <= pivot_out_2_37;
         start_in_2_38 <= start_out_2_37;
     end

     always @(posedge clk) begin
         data_in_2_38 <= data_out_1_38;
     end
  
     processor_AB AB_2_38 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_38),
       .start_in   (start_in_2_38),
       .op_in      (op_in_2_38),
       .pivot_in   (pivot_in_2_38),
       .start_out  (start_out_2_38),
       .data_out   (data_out_2_38),
       .op_out     (op_out_2_38),
       .pivot_out  (pivot_out_2_38),
       .r          (r_2_38)
     );

  // row 2, col 39

     reg start_in_2_39;
     wire start_out_2_39;

     reg [1:0] op_in_2_39;
     wire [1:0] op_out_2_39;

     wire r_2_39;

     reg data_in_2_39;
     wire data_out_2_39;

     reg pivot_in_2_39;
     wire pivot_out_2_39;

     always @(posedge clk) begin
         op_in_2_39 <= op_out_2_38;
         pivot_in_2_39 <= pivot_out_2_38;
         start_in_2_39 <= start_out_2_38;
     end

     always @(posedge clk) begin
         data_in_2_39 <= data_out_1_39;
     end
  
     processor_AB AB_2_39 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_39),
       .start_in   (start_in_2_39),
       .op_in      (op_in_2_39),
       .pivot_in   (pivot_in_2_39),
       .start_out  (start_out_2_39),
       .data_out   (data_out_2_39),
       .op_out     (op_out_2_39),
       .pivot_out  (pivot_out_2_39),
       .r          (r_2_39)
     );

  // row 2, col 40

     reg start_in_2_40;
     wire start_out_2_40;

     reg [1:0] op_in_2_40;
     wire [1:0] op_out_2_40;

     wire r_2_40;

     reg data_in_2_40;
     wire data_out_2_40;

     reg pivot_in_2_40;
     wire pivot_out_2_40;

     always @(posedge clk) begin
         op_in_2_40 <= op_out_2_39;
         pivot_in_2_40 <= pivot_out_2_39;
         start_in_2_40 <= start_out_2_39;
     end

     always @(posedge clk) begin
         data_in_2_40 <= data_out_1_40;
     end
  
     processor_AB AB_2_40 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_40),
       .start_in   (start_in_2_40),
       .op_in      (op_in_2_40),
       .pivot_in   (pivot_in_2_40),
       .start_out  (start_out_2_40),
       .data_out   (data_out_2_40),
       .op_out     (op_out_2_40),
       .pivot_out  (pivot_out_2_40),
       .r          (r_2_40)
     );

  // row 2, col 41

     reg start_in_2_41;
     wire start_out_2_41;

     reg [1:0] op_in_2_41;
     wire [1:0] op_out_2_41;

     wire r_2_41;

     reg data_in_2_41;
     wire data_out_2_41;

     reg pivot_in_2_41;
     wire pivot_out_2_41;

     always @(posedge clk) begin
         op_in_2_41 <= op_out_2_40;
         pivot_in_2_41 <= pivot_out_2_40;
         start_in_2_41 <= start_out_2_40;
     end

     always @(posedge clk) begin
         data_in_2_41 <= data_out_1_41;
     end
  
     processor_AB AB_2_41 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_41),
       .start_in   (start_in_2_41),
       .op_in      (op_in_2_41),
       .pivot_in   (pivot_in_2_41),
       .start_out  (start_out_2_41),
       .data_out   (data_out_2_41),
       .op_out     (op_out_2_41),
       .pivot_out  (pivot_out_2_41),
       .r          (r_2_41)
     );

  // row 2, col 42

     reg start_in_2_42;
     wire start_out_2_42;

     reg [1:0] op_in_2_42;
     wire [1:0] op_out_2_42;

     wire r_2_42;

     reg data_in_2_42;
     wire data_out_2_42;

     reg pivot_in_2_42;
     wire pivot_out_2_42;

     always @(posedge clk) begin
         op_in_2_42 <= op_out_2_41;
         pivot_in_2_42 <= pivot_out_2_41;
         start_in_2_42 <= start_out_2_41;
     end

     always @(posedge clk) begin
         data_in_2_42 <= data_out_1_42;
     end
  
     processor_AB AB_2_42 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_42),
       .start_in   (start_in_2_42),
       .op_in      (op_in_2_42),
       .pivot_in   (pivot_in_2_42),
       .start_out  (start_out_2_42),
       .data_out   (data_out_2_42),
       .op_out     (op_out_2_42),
       .pivot_out  (pivot_out_2_42),
       .r          (r_2_42)
     );

  // row 2, col 43

     reg start_in_2_43;
     wire start_out_2_43;

     reg [1:0] op_in_2_43;
     wire [1:0] op_out_2_43;

     wire r_2_43;

     reg data_in_2_43;
     wire data_out_2_43;

     reg pivot_in_2_43;
     wire pivot_out_2_43;

     always @(posedge clk) begin
         op_in_2_43 <= op_out_2_42;
         pivot_in_2_43 <= pivot_out_2_42;
         start_in_2_43 <= start_out_2_42;
     end

     always @(posedge clk) begin
         data_in_2_43 <= data_out_1_43;
     end
  
     processor_AB AB_2_43 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_43),
       .start_in   (start_in_2_43),
       .op_in      (op_in_2_43),
       .pivot_in   (pivot_in_2_43),
       .start_out  (start_out_2_43),
       .data_out   (data_out_2_43),
       .op_out     (op_out_2_43),
       .pivot_out  (pivot_out_2_43),
       .r          (r_2_43)
     );

  // row 2, col 44

     reg start_in_2_44;
     wire start_out_2_44;

     reg [1:0] op_in_2_44;
     wire [1:0] op_out_2_44;

     wire r_2_44;

     reg data_in_2_44;
     wire data_out_2_44;

     reg pivot_in_2_44;
     wire pivot_out_2_44;

     always @(posedge clk) begin
         op_in_2_44 <= op_out_2_43;
         pivot_in_2_44 <= pivot_out_2_43;
         start_in_2_44 <= start_out_2_43;
     end

     always @(posedge clk) begin
         data_in_2_44 <= data_out_1_44;
     end
  
     processor_AB AB_2_44 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_44),
       .start_in   (start_in_2_44),
       .op_in      (op_in_2_44),
       .pivot_in   (pivot_in_2_44),
       .start_out  (start_out_2_44),
       .data_out   (data_out_2_44),
       .op_out     (op_out_2_44),
       .pivot_out  (pivot_out_2_44),
       .r          (r_2_44)
     );

  // row 2, col 45

     reg start_in_2_45;
     wire start_out_2_45;

     reg [1:0] op_in_2_45;
     wire [1:0] op_out_2_45;

     wire r_2_45;

     reg data_in_2_45;
     wire data_out_2_45;

     reg pivot_in_2_45;
     wire pivot_out_2_45;

     always @(posedge clk) begin
         op_in_2_45 <= op_out_2_44;
         pivot_in_2_45 <= pivot_out_2_44;
         start_in_2_45 <= start_out_2_44;
     end

     always @(posedge clk) begin
         data_in_2_45 <= data_out_1_45;
     end
  
     processor_AB AB_2_45 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_45),
       .start_in   (start_in_2_45),
       .op_in      (op_in_2_45),
       .pivot_in   (pivot_in_2_45),
       .start_out  (start_out_2_45),
       .data_out   (data_out_2_45),
       .op_out     (op_out_2_45),
       .pivot_out  (pivot_out_2_45),
       .r          (r_2_45)
     );

  // row 2, col 46

     reg start_in_2_46;
     wire start_out_2_46;

     reg [1:0] op_in_2_46;
     wire [1:0] op_out_2_46;

     wire r_2_46;

     reg data_in_2_46;
     wire data_out_2_46;

     reg pivot_in_2_46;
     wire pivot_out_2_46;

     always @(posedge clk) begin
         op_in_2_46 <= op_out_2_45;
         pivot_in_2_46 <= pivot_out_2_45;
         start_in_2_46 <= start_out_2_45;
     end

     always @(posedge clk) begin
         data_in_2_46 <= data_out_1_46;
     end
  
     processor_AB AB_2_46 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_46),
       .start_in   (start_in_2_46),
       .op_in      (op_in_2_46),
       .pivot_in   (pivot_in_2_46),
       .start_out  (start_out_2_46),
       .data_out   (data_out_2_46),
       .op_out     (op_out_2_46),
       .pivot_out  (pivot_out_2_46),
       .r          (r_2_46)
     );

  // row 2, col 47

     reg start_in_2_47;
     wire start_out_2_47;

     reg [1:0] op_in_2_47;
     wire [1:0] op_out_2_47;

     wire r_2_47;

     reg data_in_2_47;
     wire data_out_2_47;

     reg pivot_in_2_47;
     wire pivot_out_2_47;

     always @(posedge clk) begin
         op_in_2_47 <= op_out_2_46;
         pivot_in_2_47 <= pivot_out_2_46;
         start_in_2_47 <= start_out_2_46;
     end

     always @(posedge clk) begin
         data_in_2_47 <= data_out_1_47;
     end
  
     processor_AB AB_2_47 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_47),
       .start_in   (start_in_2_47),
       .op_in      (op_in_2_47),
       .pivot_in   (pivot_in_2_47),
       .start_out  (start_out_2_47),
       .data_out   (data_out_2_47),
       .op_out     (op_out_2_47),
       .pivot_out  (pivot_out_2_47),
       .r          (r_2_47)
     );

  // row 2, col 48

     reg start_in_2_48;
     wire start_out_2_48;

     reg [1:0] op_in_2_48;
     wire [1:0] op_out_2_48;

     wire r_2_48;

     reg data_in_2_48;
     wire data_out_2_48;

     reg pivot_in_2_48;
     wire pivot_out_2_48;

     always @(posedge clk) begin
         op_in_2_48 <= op_out_2_47;
         pivot_in_2_48 <= pivot_out_2_47;
         start_in_2_48 <= start_out_2_47;
     end

     always @(posedge clk) begin
         data_in_2_48 <= data_out_1_48;
     end
  
     processor_AB AB_2_48 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_48),
       .start_in   (start_in_2_48),
       .op_in      (op_in_2_48),
       .pivot_in   (pivot_in_2_48),
       .start_out  (start_out_2_48),
       .data_out   (data_out_2_48),
       .op_out     (op_out_2_48),
       .pivot_out  (pivot_out_2_48),
       .r          (r_2_48)
     );

  // row 2, col 49

     reg start_in_2_49;
     wire start_out_2_49;

     reg [1:0] op_in_2_49;
     wire [1:0] op_out_2_49;

     wire r_2_49;

     reg data_in_2_49;
     wire data_out_2_49;

     reg pivot_in_2_49;
     wire pivot_out_2_49;

     always @(posedge clk) begin
         op_in_2_49 <= op_out_2_48;
         pivot_in_2_49 <= pivot_out_2_48;
         start_in_2_49 <= start_out_2_48;
     end

     always @(posedge clk) begin
         data_in_2_49 <= data_out_1_49;
     end
  
     processor_AB AB_2_49 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_49),
       .start_in   (start_in_2_49),
       .op_in      (op_in_2_49),
       .pivot_in   (pivot_in_2_49),
       .start_out  (start_out_2_49),
       .data_out   (data_out_2_49),
       .op_out     (op_out_2_49),
       .pivot_out  (pivot_out_2_49),
       .r          (r_2_49)
     );

  // row 2, col 50

     reg start_in_2_50;
     wire start_out_2_50;

     reg [1:0] op_in_2_50;
     wire [1:0] op_out_2_50;

     wire r_2_50;

     reg data_in_2_50;
     wire data_out_2_50;

     reg pivot_in_2_50;
     wire pivot_out_2_50;

     always @(posedge clk) begin
         op_in_2_50 <= op_out_2_49;
         pivot_in_2_50 <= pivot_out_2_49;
         start_in_2_50 <= start_out_2_49;
     end

     always @(posedge clk) begin
         data_in_2_50 <= data_out_1_50;
     end
  
     processor_AB AB_2_50 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_50),
       .start_in   (start_in_2_50),
       .op_in      (op_in_2_50),
       .pivot_in   (pivot_in_2_50),
       .start_out  (start_out_2_50),
       .data_out   (data_out_2_50),
       .op_out     (op_out_2_50),
       .pivot_out  (pivot_out_2_50),
       .r          (r_2_50)
     );

  // row 2, col 51

     reg start_in_2_51;
     wire start_out_2_51;

     reg [1:0] op_in_2_51;
     wire [1:0] op_out_2_51;

     wire r_2_51;

     reg data_in_2_51;
     wire data_out_2_51;

     reg pivot_in_2_51;
     wire pivot_out_2_51;

     always @(posedge clk) begin
         op_in_2_51 <= op_out_2_50;
         pivot_in_2_51 <= pivot_out_2_50;
         start_in_2_51 <= start_out_2_50;
     end

     always @(posedge clk) begin
         data_in_2_51 <= data_out_1_51;
     end
  
     processor_AB AB_2_51 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_51),
       .start_in   (start_in_2_51),
       .op_in      (op_in_2_51),
       .pivot_in   (pivot_in_2_51),
       .start_out  (start_out_2_51),
       .data_out   (data_out_2_51),
       .op_out     (op_out_2_51),
       .pivot_out  (pivot_out_2_51),
       .r          (r_2_51)
     );

  // row 2, col 52

     reg start_in_2_52;
     wire start_out_2_52;

     reg [1:0] op_in_2_52;
     wire [1:0] op_out_2_52;

     wire r_2_52;

     reg data_in_2_52;
     wire data_out_2_52;

     reg pivot_in_2_52;
     wire pivot_out_2_52;

     always @(posedge clk) begin
         op_in_2_52 <= op_out_2_51;
         pivot_in_2_52 <= pivot_out_2_51;
         start_in_2_52 <= start_out_2_51;
     end

     always @(posedge clk) begin
         data_in_2_52 <= data_out_1_52;
     end
  
     processor_AB AB_2_52 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_52),
       .start_in   (start_in_2_52),
       .op_in      (op_in_2_52),
       .pivot_in   (pivot_in_2_52),
       .start_out  (start_out_2_52),
       .data_out   (data_out_2_52),
       .op_out     (op_out_2_52),
       .pivot_out  (pivot_out_2_52),
       .r          (r_2_52)
     );

  // row 2, col 53

     reg start_in_2_53;
     wire start_out_2_53;

     reg [1:0] op_in_2_53;
     wire [1:0] op_out_2_53;

     wire r_2_53;

     reg data_in_2_53;
     wire data_out_2_53;

     reg pivot_in_2_53;
     wire pivot_out_2_53;

     always @(posedge clk) begin
         op_in_2_53 <= op_out_2_52;
         pivot_in_2_53 <= pivot_out_2_52;
         start_in_2_53 <= start_out_2_52;
     end

     always @(posedge clk) begin
         data_in_2_53 <= data_out_1_53;
     end
  
     processor_AB AB_2_53 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_53),
       .start_in   (start_in_2_53),
       .op_in      (op_in_2_53),
       .pivot_in   (pivot_in_2_53),
       .start_out  (start_out_2_53),
       .data_out   (data_out_2_53),
       .op_out     (op_out_2_53),
       .pivot_out  (pivot_out_2_53),
       .r          (r_2_53)
     );

  // row 2, col 54

     reg start_in_2_54;
     wire start_out_2_54;

     reg [1:0] op_in_2_54;
     wire [1:0] op_out_2_54;

     wire r_2_54;

     reg data_in_2_54;
     wire data_out_2_54;

     reg pivot_in_2_54;
     wire pivot_out_2_54;

     always @(posedge clk) begin
         op_in_2_54 <= op_out_2_53;
         pivot_in_2_54 <= pivot_out_2_53;
         start_in_2_54 <= start_out_2_53;
     end

     always @(posedge clk) begin
         data_in_2_54 <= data_out_1_54;
     end
  
     processor_AB AB_2_54 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_54),
       .start_in   (start_in_2_54),
       .op_in      (op_in_2_54),
       .pivot_in   (pivot_in_2_54),
       .start_out  (start_out_2_54),
       .data_out   (data_out_2_54),
       .op_out     (op_out_2_54),
       .pivot_out  (pivot_out_2_54),
       .r          (r_2_54)
     );

  // row 2, col 55

     reg start_in_2_55;
     wire start_out_2_55;

     reg [1:0] op_in_2_55;
     wire [1:0] op_out_2_55;

     wire r_2_55;

     reg data_in_2_55;
     wire data_out_2_55;

     reg pivot_in_2_55;
     wire pivot_out_2_55;

     always @(posedge clk) begin
         op_in_2_55 <= op_out_2_54;
         pivot_in_2_55 <= pivot_out_2_54;
         start_in_2_55 <= start_out_2_54;
     end

     always @(posedge clk) begin
         data_in_2_55 <= data_out_1_55;
     end
  
     processor_AB AB_2_55 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_55),
       .start_in   (start_in_2_55),
       .op_in      (op_in_2_55),
       .pivot_in   (pivot_in_2_55),
       .start_out  (start_out_2_55),
       .data_out   (data_out_2_55),
       .op_out     (op_out_2_55),
       .pivot_out  (pivot_out_2_55),
       .r          (r_2_55)
     );

  // row 2, col 56

     reg start_in_2_56;
     wire start_out_2_56;

     reg [1:0] op_in_2_56;
     wire [1:0] op_out_2_56;

     wire r_2_56;

     reg data_in_2_56;
     wire data_out_2_56;

     reg pivot_in_2_56;
     wire pivot_out_2_56;

     always @(posedge clk) begin
         op_in_2_56 <= op_out_2_55;
         pivot_in_2_56 <= pivot_out_2_55;
         start_in_2_56 <= start_out_2_55;
     end

     always @(posedge clk) begin
         data_in_2_56 <= data_out_1_56;
     end
  
     processor_AB AB_2_56 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_56),
       .start_in   (start_in_2_56),
       .op_in      (op_in_2_56),
       .pivot_in   (pivot_in_2_56),
       .start_out  (start_out_2_56),
       .data_out   (data_out_2_56),
       .op_out     (op_out_2_56),
       .pivot_out  (pivot_out_2_56),
       .r          (r_2_56)
     );

  // row 2, col 57

     reg start_in_2_57;
     wire start_out_2_57;

     reg [1:0] op_in_2_57;
     wire [1:0] op_out_2_57;

     wire r_2_57;

     reg data_in_2_57;
     wire data_out_2_57;

     reg pivot_in_2_57;
     wire pivot_out_2_57;

     always @(posedge clk) begin
         op_in_2_57 <= op_out_2_56;
         pivot_in_2_57 <= pivot_out_2_56;
         start_in_2_57 <= start_out_2_56;
     end

     always @(posedge clk) begin
         data_in_2_57 <= data_out_1_57;
     end
  
     processor_AB AB_2_57 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_57),
       .start_in   (start_in_2_57),
       .op_in      (op_in_2_57),
       .pivot_in   (pivot_in_2_57),
       .start_out  (start_out_2_57),
       .data_out   (data_out_2_57),
       .op_out     (op_out_2_57),
       .pivot_out  (pivot_out_2_57),
       .r          (r_2_57)
     );

  // row 2, col 58

     reg start_in_2_58;
     wire start_out_2_58;

     reg [1:0] op_in_2_58;
     wire [1:0] op_out_2_58;

     wire r_2_58;

     reg data_in_2_58;
     wire data_out_2_58;

     reg pivot_in_2_58;
     wire pivot_out_2_58;

     always @(posedge clk) begin
         op_in_2_58 <= op_out_2_57;
         pivot_in_2_58 <= pivot_out_2_57;
         start_in_2_58 <= start_out_2_57;
     end

     always @(posedge clk) begin
         data_in_2_58 <= data_out_1_58;
     end
  
     processor_AB AB_2_58 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_58),
       .start_in   (start_in_2_58),
       .op_in      (op_in_2_58),
       .pivot_in   (pivot_in_2_58),
       .start_out  (start_out_2_58),
       .data_out   (data_out_2_58),
       .op_out     (op_out_2_58),
       .pivot_out  (pivot_out_2_58),
       .r          (r_2_58)
     );

  // row 2, col 59

     reg start_in_2_59;
     wire start_out_2_59;

     reg [1:0] op_in_2_59;
     wire [1:0] op_out_2_59;

     wire r_2_59;

     reg data_in_2_59;
     wire data_out_2_59;

     reg pivot_in_2_59;
     wire pivot_out_2_59;

     always @(posedge clk) begin
         op_in_2_59 <= op_out_2_58;
         pivot_in_2_59 <= pivot_out_2_58;
         start_in_2_59 <= start_out_2_58;
     end

     always @(posedge clk) begin
         data_in_2_59 <= data_out_1_59;
     end
  
     processor_AB AB_2_59 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_59),
       .start_in   (start_in_2_59),
       .op_in      (op_in_2_59),
       .pivot_in   (pivot_in_2_59),
       .start_out  (start_out_2_59),
       .data_out   (data_out_2_59),
       .op_out     (op_out_2_59),
       .pivot_out  (pivot_out_2_59),
       .r          (r_2_59)
     );

  // row 2, col 60

     reg start_in_2_60;
     wire start_out_2_60;

     reg [1:0] op_in_2_60;
     wire [1:0] op_out_2_60;

     wire r_2_60;

     reg data_in_2_60;
     wire data_out_2_60;

     reg pivot_in_2_60;
     wire pivot_out_2_60;

     always @(posedge clk) begin
         op_in_2_60 <= op_out_2_59;
         pivot_in_2_60 <= pivot_out_2_59;
         start_in_2_60 <= start_out_2_59;
     end

     always @(posedge clk) begin
         data_in_2_60 <= data_out_1_60;
     end
  
     processor_AB AB_2_60 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_60),
       .start_in   (start_in_2_60),
       .op_in      (op_in_2_60),
       .pivot_in   (pivot_in_2_60),
       .start_out  (start_out_2_60),
       .data_out   (data_out_2_60),
       .op_out     (op_out_2_60),
       .pivot_out  (pivot_out_2_60),
       .r          (r_2_60)
     );

  // row 2, col 61

     reg start_in_2_61;
     wire start_out_2_61;

     reg [1:0] op_in_2_61;
     wire [1:0] op_out_2_61;

     wire r_2_61;

     reg data_in_2_61;
     wire data_out_2_61;

     reg pivot_in_2_61;
     wire pivot_out_2_61;

     always @(posedge clk) begin
         op_in_2_61 <= op_out_2_60;
         pivot_in_2_61 <= pivot_out_2_60;
         start_in_2_61 <= start_out_2_60;
     end

     always @(posedge clk) begin
         data_in_2_61 <= data_out_1_61;
     end
  
     processor_AB AB_2_61 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_61),
       .start_in   (start_in_2_61),
       .op_in      (op_in_2_61),
       .pivot_in   (pivot_in_2_61),
       .start_out  (start_out_2_61),
       .data_out   (data_out_2_61),
       .op_out     (op_out_2_61),
       .pivot_out  (pivot_out_2_61),
       .r          (r_2_61)
     );

  // row 2, col 62

     reg start_in_2_62;
     wire start_out_2_62;

     reg [1:0] op_in_2_62;
     wire [1:0] op_out_2_62;

     wire r_2_62;

     reg data_in_2_62;
     wire data_out_2_62;

     reg pivot_in_2_62;
     wire pivot_out_2_62;

     always @(posedge clk) begin
         op_in_2_62 <= op_out_2_61;
         pivot_in_2_62 <= pivot_out_2_61;
         start_in_2_62 <= start_out_2_61;
     end

     always @(posedge clk) begin
         data_in_2_62 <= data_out_1_62;
     end
  
     processor_AB AB_2_62 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_62),
       .start_in   (start_in_2_62),
       .op_in      (op_in_2_62),
       .pivot_in   (pivot_in_2_62),
       .start_out  (start_out_2_62),
       .data_out   (data_out_2_62),
       .op_out     (op_out_2_62),
       .pivot_out  (pivot_out_2_62),
       .r          (r_2_62)
     );

  // row 2, col 63

     reg start_in_2_63;
     wire start_out_2_63;

     reg [1:0] op_in_2_63;
     wire [1:0] op_out_2_63;

     wire r_2_63;

     reg data_in_2_63;
     wire data_out_2_63;

     reg pivot_in_2_63;
     wire pivot_out_2_63;

     always @(posedge clk) begin
         op_in_2_63 <= op_out_2_62;
         pivot_in_2_63 <= pivot_out_2_62;
         start_in_2_63 <= start_out_2_62;
     end

     always @(posedge clk) begin
         data_in_2_63 <= data_out_1_63;
     end
  
     processor_AB AB_2_63 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_63),
       .start_in   (start_in_2_63),
       .op_in      (op_in_2_63),
       .pivot_in   (pivot_in_2_63),
       .start_out  (start_out_2_63),
       .data_out   (data_out_2_63),
       .op_out     (op_out_2_63),
       .pivot_out  (pivot_out_2_63),
       .r          (r_2_63)
     );

  // row 2, col 64

     reg start_in_2_64;
     wire start_out_2_64;

     reg [1:0] op_in_2_64;
     wire [1:0] op_out_2_64;

     wire r_2_64;

     reg data_in_2_64;
     wire data_out_2_64;

     reg pivot_in_2_64;
     wire pivot_out_2_64;

     always @(posedge clk) begin
         op_in_2_64 <= op_out_2_63;
         pivot_in_2_64 <= pivot_out_2_63;
         start_in_2_64 <= start_out_2_63;
     end

     always @(posedge clk) begin
         data_in_2_64 <= data_out_1_64;
     end
  
     processor_AB AB_2_64 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_64),
       .start_in   (start_in_2_64),
       .op_in      (op_in_2_64),
       .pivot_in   (pivot_in_2_64),
       .start_out  (start_out_2_64),
       .data_out   (data_out_2_64),
       .op_out     (op_out_2_64),
       .pivot_out  (pivot_out_2_64),
       .r          (r_2_64)
     );

  // row 2, col 65

     reg start_in_2_65;
     wire start_out_2_65;

     reg [1:0] op_in_2_65;
     wire [1:0] op_out_2_65;

     wire r_2_65;

     reg data_in_2_65;
     wire data_out_2_65;

     reg pivot_in_2_65;
     wire pivot_out_2_65;

     always @(posedge clk) begin
         op_in_2_65 <= op_out_2_64;
         pivot_in_2_65 <= pivot_out_2_64;
         start_in_2_65 <= start_out_2_64;
     end

     always @(posedge clk) begin
         data_in_2_65 <= data_out_1_65;
     end
  
     processor_AB AB_2_65 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_65),
       .start_in   (start_in_2_65),
       .op_in      (op_in_2_65),
       .pivot_in   (pivot_in_2_65),
       .start_out  (start_out_2_65),
       .data_out   (data_out_2_65),
       .op_out     (op_out_2_65),
       .pivot_out  (pivot_out_2_65),
       .r          (r_2_65)
     );

  // row 2, col 66

     reg start_in_2_66;
     wire start_out_2_66;

     reg [1:0] op_in_2_66;
     wire [1:0] op_out_2_66;

     wire r_2_66;

     reg data_in_2_66;
     wire data_out_2_66;

     reg pivot_in_2_66;
     wire pivot_out_2_66;

     always @(posedge clk) begin
         op_in_2_66 <= op_out_2_65;
         pivot_in_2_66 <= pivot_out_2_65;
         start_in_2_66 <= start_out_2_65;
     end

     always @(posedge clk) begin
         data_in_2_66 <= data_out_1_66;
     end
  
     processor_AB AB_2_66 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_66),
       .start_in   (start_in_2_66),
       .op_in      (op_in_2_66),
       .pivot_in   (pivot_in_2_66),
       .start_out  (start_out_2_66),
       .data_out   (data_out_2_66),
       .op_out     (op_out_2_66),
       .pivot_out  (pivot_out_2_66),
       .r          (r_2_66)
     );

  // row 2, col 67

     reg start_in_2_67;
     wire start_out_2_67;

     reg [1:0] op_in_2_67;
     wire [1:0] op_out_2_67;

     wire r_2_67;

     reg data_in_2_67;
     wire data_out_2_67;

     reg pivot_in_2_67;
     wire pivot_out_2_67;

     always @(posedge clk) begin
         op_in_2_67 <= op_out_2_66;
         pivot_in_2_67 <= pivot_out_2_66;
         start_in_2_67 <= start_out_2_66;
     end

     always @(posedge clk) begin
         data_in_2_67 <= data_out_1_67;
     end
  
     processor_AB AB_2_67 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_67),
       .start_in   (start_in_2_67),
       .op_in      (op_in_2_67),
       .pivot_in   (pivot_in_2_67),
       .start_out  (start_out_2_67),
       .data_out   (data_out_2_67),
       .op_out     (op_out_2_67),
       .pivot_out  (pivot_out_2_67),
       .r          (r_2_67)
     );

  // row 2, col 68

     reg start_in_2_68;
     wire start_out_2_68;

     reg [1:0] op_in_2_68;
     wire [1:0] op_out_2_68;

     wire r_2_68;

     reg data_in_2_68;
     wire data_out_2_68;

     reg pivot_in_2_68;
     wire pivot_out_2_68;

     always @(posedge clk) begin
         op_in_2_68 <= op_out_2_67;
         pivot_in_2_68 <= pivot_out_2_67;
         start_in_2_68 <= start_out_2_67;
     end

     always @(posedge clk) begin
         data_in_2_68 <= data_out_1_68;
     end
  
     processor_AB AB_2_68 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_68),
       .start_in   (start_in_2_68),
       .op_in      (op_in_2_68),
       .pivot_in   (pivot_in_2_68),
       .start_out  (start_out_2_68),
       .data_out   (data_out_2_68),
       .op_out     (op_out_2_68),
       .pivot_out  (pivot_out_2_68),
       .r          (r_2_68)
     );

  // row 2, col 69

     reg start_in_2_69;
     wire start_out_2_69;

     reg [1:0] op_in_2_69;
     wire [1:0] op_out_2_69;

     wire r_2_69;

     reg data_in_2_69;
     wire data_out_2_69;

     reg pivot_in_2_69;
     wire pivot_out_2_69;

     always @(posedge clk) begin
         op_in_2_69 <= op_out_2_68;
         pivot_in_2_69 <= pivot_out_2_68;
         start_in_2_69 <= start_out_2_68;
     end

     always @(posedge clk) begin
         data_in_2_69 <= data_out_1_69;
     end
  
     processor_AB AB_2_69 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_69),
       .start_in   (start_in_2_69),
       .op_in      (op_in_2_69),
       .pivot_in   (pivot_in_2_69),
       .start_out  (start_out_2_69),
       .data_out   (data_out_2_69),
       .op_out     (op_out_2_69),
       .pivot_out  (pivot_out_2_69),
       .r          (r_2_69)
     );

  // row 2, col 70

     reg start_in_2_70;
     wire start_out_2_70;

     reg [1:0] op_in_2_70;
     wire [1:0] op_out_2_70;

     wire r_2_70;

     reg data_in_2_70;
     wire data_out_2_70;

     reg pivot_in_2_70;
     wire pivot_out_2_70;

     always @(posedge clk) begin
         op_in_2_70 <= op_out_2_69;
         pivot_in_2_70 <= pivot_out_2_69;
         start_in_2_70 <= start_out_2_69;
     end

     always @(posedge clk) begin
         data_in_2_70 <= data_out_1_70;
     end
  
     processor_AB AB_2_70 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_70),
       .start_in   (start_in_2_70),
       .op_in      (op_in_2_70),
       .pivot_in   (pivot_in_2_70),
       .start_out  (start_out_2_70),
       .data_out   (data_out_2_70),
       .op_out     (op_out_2_70),
       .pivot_out  (pivot_out_2_70),
       .r          (r_2_70)
     );

  // row 2, col 71

     reg start_in_2_71;
     wire start_out_2_71;

     reg [1:0] op_in_2_71;
     wire [1:0] op_out_2_71;

     wire r_2_71;

     reg data_in_2_71;
     wire data_out_2_71;

     reg pivot_in_2_71;
     wire pivot_out_2_71;

     always @(posedge clk) begin
         op_in_2_71 <= op_out_2_70;
         pivot_in_2_71 <= pivot_out_2_70;
         start_in_2_71 <= start_out_2_70;
     end

     always @(posedge clk) begin
         data_in_2_71 <= data_out_1_71;
     end
  
     processor_AB AB_2_71 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_71),
       .start_in   (start_in_2_71),
       .op_in      (op_in_2_71),
       .pivot_in   (pivot_in_2_71),
       .start_out  (start_out_2_71),
       .data_out   (data_out_2_71),
       .op_out     (op_out_2_71),
       .pivot_out  (pivot_out_2_71),
       .r          (r_2_71)
     );

  // row 2, col 72

     reg start_in_2_72;
     wire start_out_2_72;

     reg [1:0] op_in_2_72;
     wire [1:0] op_out_2_72;

     wire r_2_72;

     reg data_in_2_72;
     wire data_out_2_72;

     reg pivot_in_2_72;
     wire pivot_out_2_72;

     always @(posedge clk) begin
         op_in_2_72 <= op_out_2_71;
         pivot_in_2_72 <= pivot_out_2_71;
         start_in_2_72 <= start_out_2_71;
     end

     always @(posedge clk) begin
         data_in_2_72 <= data_out_1_72;
     end
  
     processor_AB AB_2_72 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_72),
       .start_in   (start_in_2_72),
       .op_in      (op_in_2_72),
       .pivot_in   (pivot_in_2_72),
       .start_out  (start_out_2_72),
       .data_out   (data_out_2_72),
       .op_out     (op_out_2_72),
       .pivot_out  (pivot_out_2_72),
       .r          (r_2_72)
     );

  // row 2, col 73

     reg start_in_2_73;
     wire start_out_2_73;

     reg [1:0] op_in_2_73;
     wire [1:0] op_out_2_73;

     wire r_2_73;

     reg data_in_2_73;
     wire data_out_2_73;

     reg pivot_in_2_73;
     wire pivot_out_2_73;

     always @(posedge clk) begin
         op_in_2_73 <= op_out_2_72;
         pivot_in_2_73 <= pivot_out_2_72;
         start_in_2_73 <= start_out_2_72;
     end

     always @(posedge clk) begin
         data_in_2_73 <= data_out_1_73;
     end
  
     processor_AB AB_2_73 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_73),
       .start_in   (start_in_2_73),
       .op_in      (op_in_2_73),
       .pivot_in   (pivot_in_2_73),
       .start_out  (start_out_2_73),
       .data_out   (data_out_2_73),
       .op_out     (op_out_2_73),
       .pivot_out  (pivot_out_2_73),
       .r          (r_2_73)
     );

  // row 2, col 74

     reg start_in_2_74;
     wire start_out_2_74;

     reg [1:0] op_in_2_74;
     wire [1:0] op_out_2_74;

     wire r_2_74;

     reg data_in_2_74;
     wire data_out_2_74;

     reg pivot_in_2_74;
     wire pivot_out_2_74;

     always @(posedge clk) begin
         op_in_2_74 <= op_out_2_73;
         pivot_in_2_74 <= pivot_out_2_73;
         start_in_2_74 <= start_out_2_73;
     end

     always @(posedge clk) begin
         data_in_2_74 <= data_out_1_74;
     end
  
     processor_AB AB_2_74 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_74),
       .start_in   (start_in_2_74),
       .op_in      (op_in_2_74),
       .pivot_in   (pivot_in_2_74),
       .start_out  (start_out_2_74),
       .data_out   (data_out_2_74),
       .op_out     (op_out_2_74),
       .pivot_out  (pivot_out_2_74),
       .r          (r_2_74)
     );

  // row 2, col 75

     reg start_in_2_75;
     wire start_out_2_75;

     reg [1:0] op_in_2_75;
     wire [1:0] op_out_2_75;

     wire r_2_75;

     reg data_in_2_75;
     wire data_out_2_75;

     reg pivot_in_2_75;
     wire pivot_out_2_75;

     always @(posedge clk) begin
         op_in_2_75 <= op_out_2_74;
         pivot_in_2_75 <= pivot_out_2_74;
         start_in_2_75 <= start_out_2_74;
     end

     always @(posedge clk) begin
         data_in_2_75 <= data_out_1_75;
     end
  
     processor_AB AB_2_75 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_75),
       .start_in   (start_in_2_75),
       .op_in      (op_in_2_75),
       .pivot_in   (pivot_in_2_75),
       .start_out  (start_out_2_75),
       .data_out   (data_out_2_75),
       .op_out     (op_out_2_75),
       .pivot_out  (pivot_out_2_75),
       .r          (r_2_75)
     );

  // row 2, col 76

     reg start_in_2_76;
     wire start_out_2_76;

     reg [1:0] op_in_2_76;
     wire [1:0] op_out_2_76;

     wire r_2_76;

     reg data_in_2_76;
     wire data_out_2_76;

     reg pivot_in_2_76;
     wire pivot_out_2_76;

     always @(posedge clk) begin
         op_in_2_76 <= op_out_2_75;
         pivot_in_2_76 <= pivot_out_2_75;
         start_in_2_76 <= start_out_2_75;
     end

     always @(posedge clk) begin
         data_in_2_76 <= data_out_1_76;
     end
  
     processor_AB AB_2_76 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_76),
       .start_in   (start_in_2_76),
       .op_in      (op_in_2_76),
       .pivot_in   (pivot_in_2_76),
       .start_out  (start_out_2_76),
       .data_out   (data_out_2_76),
       .op_out     (op_out_2_76),
       .pivot_out  (pivot_out_2_76),
       .r          (r_2_76)
     );

  // row 2, col 77

     reg start_in_2_77;
     wire start_out_2_77;

     reg [1:0] op_in_2_77;
     wire [1:0] op_out_2_77;

     wire r_2_77;

     reg data_in_2_77;
     wire data_out_2_77;

     reg pivot_in_2_77;
     wire pivot_out_2_77;

     always @(posedge clk) begin
         op_in_2_77 <= op_out_2_76;
         pivot_in_2_77 <= pivot_out_2_76;
         start_in_2_77 <= start_out_2_76;
     end

     always @(posedge clk) begin
         data_in_2_77 <= data_out_1_77;
     end
  
     processor_AB AB_2_77 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_77),
       .start_in   (start_in_2_77),
       .op_in      (op_in_2_77),
       .pivot_in   (pivot_in_2_77),
       .start_out  (start_out_2_77),
       .data_out   (data_out_2_77),
       .op_out     (op_out_2_77),
       .pivot_out  (pivot_out_2_77),
       .r          (r_2_77)
     );

  // row 2, col 78

     reg start_in_2_78;
     wire start_out_2_78;

     reg [1:0] op_in_2_78;
     wire [1:0] op_out_2_78;

     wire r_2_78;

     reg data_in_2_78;
     wire data_out_2_78;

     reg pivot_in_2_78;
     wire pivot_out_2_78;

     always @(posedge clk) begin
         op_in_2_78 <= op_out_2_77;
         pivot_in_2_78 <= pivot_out_2_77;
         start_in_2_78 <= start_out_2_77;
     end

     always @(posedge clk) begin
         data_in_2_78 <= data_out_1_78;
     end
  
     processor_AB AB_2_78 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_78),
       .start_in   (start_in_2_78),
       .op_in      (op_in_2_78),
       .pivot_in   (pivot_in_2_78),
       .start_out  (start_out_2_78),
       .data_out   (data_out_2_78),
       .op_out     (op_out_2_78),
       .pivot_out  (pivot_out_2_78),
       .r          (r_2_78)
     );

  // row 2, col 79

     reg start_in_2_79;
     wire start_out_2_79;

     reg [1:0] op_in_2_79;
     wire [1:0] op_out_2_79;

     wire r_2_79;

     reg data_in_2_79;
     wire data_out_2_79;

     reg pivot_in_2_79;
     wire pivot_out_2_79;

     always @(posedge clk) begin
         op_in_2_79 <= op_out_2_78;
         pivot_in_2_79 <= pivot_out_2_78;
         start_in_2_79 <= start_out_2_78;
     end

     always @(posedge clk) begin
         data_in_2_79 <= data_out_1_79;
     end
  
     processor_AB AB_2_79 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_79),
       .start_in   (start_in_2_79),
       .op_in      (op_in_2_79),
       .pivot_in   (pivot_in_2_79),
       .start_out  (start_out_2_79),
       .data_out   (data_out_2_79),
       .op_out     (op_out_2_79),
       .pivot_out  (pivot_out_2_79),
       .r          (r_2_79)
     );

  // row 2, col 80

     reg start_in_2_80;
     wire start_out_2_80;

     reg [1:0] op_in_2_80;
     wire [1:0] op_out_2_80;

     wire r_2_80;

     reg data_in_2_80;
     wire data_out_2_80;

     reg pivot_in_2_80;
     wire pivot_out_2_80;

     always @(posedge clk) begin
         op_in_2_80 <= op_out_2_79;
         pivot_in_2_80 <= pivot_out_2_79;
         start_in_2_80 <= start_out_2_79;
     end

     always @(posedge clk) begin
         data_in_2_80 <= data_out_1_80;
     end
  
     processor_AB AB_2_80 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_80),
       .start_in   (start_in_2_80),
       .op_in      (op_in_2_80),
       .pivot_in   (pivot_in_2_80),
       .start_out  (start_out_2_80),
       .data_out   (data_out_2_80),
       .op_out     (op_out_2_80),
       .pivot_out  (pivot_out_2_80),
       .r          (r_2_80)
     );

  // row 2, col 81

     reg start_in_2_81;
     wire start_out_2_81;

     reg [1:0] op_in_2_81;
     wire [1:0] op_out_2_81;

     wire r_2_81;

     reg data_in_2_81;
     wire data_out_2_81;

     reg pivot_in_2_81;
     wire pivot_out_2_81;

     always @(posedge clk) begin
         op_in_2_81 <= op_out_2_80;
         pivot_in_2_81 <= pivot_out_2_80;
         start_in_2_81 <= start_out_2_80;
     end

     always @(posedge clk) begin
         data_in_2_81 <= data_out_1_81;
     end
  
     processor_AB AB_2_81 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_81),
       .start_in   (start_in_2_81),
       .op_in      (op_in_2_81),
       .pivot_in   (pivot_in_2_81),
       .start_out  (start_out_2_81),
       .data_out   (data_out_2_81),
       .op_out     (op_out_2_81),
       .pivot_out  (pivot_out_2_81),
       .r          (r_2_81)
     );

  // row 2, col 82

     reg start_in_2_82;
     wire start_out_2_82;

     reg [1:0] op_in_2_82;
     wire [1:0] op_out_2_82;

     wire r_2_82;

     reg data_in_2_82;
     wire data_out_2_82;

     reg pivot_in_2_82;
     wire pivot_out_2_82;

     always @(posedge clk) begin
         op_in_2_82 <= op_out_2_81;
         pivot_in_2_82 <= pivot_out_2_81;
         start_in_2_82 <= start_out_2_81;
     end

     always @(posedge clk) begin
         data_in_2_82 <= data_out_1_82;
     end
  
     processor_AB AB_2_82 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_82),
       .start_in   (start_in_2_82),
       .op_in      (op_in_2_82),
       .pivot_in   (pivot_in_2_82),
       .start_out  (start_out_2_82),
       .data_out   (data_out_2_82),
       .op_out     (op_out_2_82),
       .pivot_out  (pivot_out_2_82),
       .r          (r_2_82)
     );

  // row 2, col 83

     reg start_in_2_83;
     wire start_out_2_83;

     reg [1:0] op_in_2_83;
     wire [1:0] op_out_2_83;

     wire r_2_83;

     reg data_in_2_83;
     wire data_out_2_83;

     reg pivot_in_2_83;
     wire pivot_out_2_83;

     always @(posedge clk) begin
         op_in_2_83 <= op_out_2_82;
         pivot_in_2_83 <= pivot_out_2_82;
         start_in_2_83 <= start_out_2_82;
     end

     always @(posedge clk) begin
         data_in_2_83 <= data_out_1_83;
     end
  
     processor_AB AB_2_83 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_83),
       .start_in   (start_in_2_83),
       .op_in      (op_in_2_83),
       .pivot_in   (pivot_in_2_83),
       .start_out  (start_out_2_83),
       .data_out   (data_out_2_83),
       .op_out     (op_out_2_83),
       .pivot_out  (pivot_out_2_83),
       .r          (r_2_83)
     );

  // row 2, col 84

     reg start_in_2_84;
     wire start_out_2_84;

     reg [1:0] op_in_2_84;
     wire [1:0] op_out_2_84;

     wire r_2_84;

     reg data_in_2_84;
     wire data_out_2_84;

     reg pivot_in_2_84;
     wire pivot_out_2_84;

     always @(posedge clk) begin
         op_in_2_84 <= op_out_2_83;
         pivot_in_2_84 <= pivot_out_2_83;
         start_in_2_84 <= start_out_2_83;
     end

     always @(posedge clk) begin
         data_in_2_84 <= data_out_1_84;
     end
  
     processor_AB AB_2_84 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_84),
       .start_in   (start_in_2_84),
       .op_in      (op_in_2_84),
       .pivot_in   (pivot_in_2_84),
       .start_out  (start_out_2_84),
       .data_out   (data_out_2_84),
       .op_out     (op_out_2_84),
       .pivot_out  (pivot_out_2_84),
       .r          (r_2_84)
     );

  // row 2, col 85

     reg start_in_2_85;
     wire start_out_2_85;

     reg [1:0] op_in_2_85;
     wire [1:0] op_out_2_85;

     wire r_2_85;

     reg data_in_2_85;
     wire data_out_2_85;

     reg pivot_in_2_85;
     wire pivot_out_2_85;

     always @(posedge clk) begin
         op_in_2_85 <= op_out_2_84;
         pivot_in_2_85 <= pivot_out_2_84;
         start_in_2_85 <= start_out_2_84;
     end

     always @(posedge clk) begin
         data_in_2_85 <= data_out_1_85;
     end
  
     processor_AB AB_2_85 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_85),
       .start_in   (start_in_2_85),
       .op_in      (op_in_2_85),
       .pivot_in   (pivot_in_2_85),
       .start_out  (start_out_2_85),
       .data_out   (data_out_2_85),
       .op_out     (op_out_2_85),
       .pivot_out  (pivot_out_2_85),
       .r          (r_2_85)
     );

  // row 2, col 86

     reg start_in_2_86;
     wire start_out_2_86;

     reg [1:0] op_in_2_86;
     wire [1:0] op_out_2_86;

     wire r_2_86;

     reg data_in_2_86;
     wire data_out_2_86;

     reg pivot_in_2_86;
     wire pivot_out_2_86;

     always @(posedge clk) begin
         op_in_2_86 <= op_out_2_85;
         pivot_in_2_86 <= pivot_out_2_85;
         start_in_2_86 <= start_out_2_85;
     end

     always @(posedge clk) begin
         data_in_2_86 <= data_out_1_86;
     end
  
     processor_AB AB_2_86 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_86),
       .start_in   (start_in_2_86),
       .op_in      (op_in_2_86),
       .pivot_in   (pivot_in_2_86),
       .start_out  (start_out_2_86),
       .data_out   (data_out_2_86),
       .op_out     (op_out_2_86),
       .pivot_out  (pivot_out_2_86),
       .r          (r_2_86)
     );

  // row 2, col 87

     reg start_in_2_87;
     wire start_out_2_87;

     reg [1:0] op_in_2_87;
     wire [1:0] op_out_2_87;

     wire r_2_87;

     reg data_in_2_87;
     wire data_out_2_87;

     reg pivot_in_2_87;
     wire pivot_out_2_87;

     always @(posedge clk) begin
         op_in_2_87 <= op_out_2_86;
         pivot_in_2_87 <= pivot_out_2_86;
         start_in_2_87 <= start_out_2_86;
     end

     always @(posedge clk) begin
         data_in_2_87 <= data_out_1_87;
     end
  
     processor_AB AB_2_87 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_87),
       .start_in   (start_in_2_87),
       .op_in      (op_in_2_87),
       .pivot_in   (pivot_in_2_87),
       .start_out  (start_out_2_87),
       .data_out   (data_out_2_87),
       .op_out     (op_out_2_87),
       .pivot_out  (pivot_out_2_87),
       .r          (r_2_87)
     );

  // row 2, col 88

     reg start_in_2_88;
     wire start_out_2_88;

     reg [1:0] op_in_2_88;
     wire [1:0] op_out_2_88;

     wire r_2_88;

     reg data_in_2_88;
     wire data_out_2_88;

     reg pivot_in_2_88;
     wire pivot_out_2_88;

     always @(posedge clk) begin
         op_in_2_88 <= op_out_2_87;
         pivot_in_2_88 <= pivot_out_2_87;
         start_in_2_88 <= start_out_2_87;
     end

     always @(posedge clk) begin
         data_in_2_88 <= data_out_1_88;
     end
  
     processor_AB AB_2_88 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_88),
       .start_in   (start_in_2_88),
       .op_in      (op_in_2_88),
       .pivot_in   (pivot_in_2_88),
       .start_out  (start_out_2_88),
       .data_out   (data_out_2_88),
       .op_out     (op_out_2_88),
       .pivot_out  (pivot_out_2_88),
       .r          (r_2_88)
     );

  // row 2, col 89

     reg start_in_2_89;
     wire start_out_2_89;

     reg [1:0] op_in_2_89;
     wire [1:0] op_out_2_89;

     wire r_2_89;

     reg data_in_2_89;
     wire data_out_2_89;

     reg pivot_in_2_89;
     wire pivot_out_2_89;

     always @(posedge clk) begin
         op_in_2_89 <= op_out_2_88;
         pivot_in_2_89 <= pivot_out_2_88;
         start_in_2_89 <= start_out_2_88;
     end

     always @(posedge clk) begin
         data_in_2_89 <= data_out_1_89;
     end
  
     processor_AB AB_2_89 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_89),
       .start_in   (start_in_2_89),
       .op_in      (op_in_2_89),
       .pivot_in   (pivot_in_2_89),
       .start_out  (start_out_2_89),
       .data_out   (data_out_2_89),
       .op_out     (op_out_2_89),
       .pivot_out  (pivot_out_2_89),
       .r          (r_2_89)
     );

  // row 2, col 90

     reg start_in_2_90;
     wire start_out_2_90;

     reg [1:0] op_in_2_90;
     wire [1:0] op_out_2_90;

     wire r_2_90;

     reg data_in_2_90;
     wire data_out_2_90;

     reg pivot_in_2_90;
     wire pivot_out_2_90;

     always @(posedge clk) begin
         op_in_2_90 <= op_out_2_89;
         pivot_in_2_90 <= pivot_out_2_89;
         start_in_2_90 <= start_out_2_89;
     end

     always @(posedge clk) begin
         data_in_2_90 <= data_out_1_90;
     end
  
     processor_AB AB_2_90 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_90),
       .start_in   (start_in_2_90),
       .op_in      (op_in_2_90),
       .pivot_in   (pivot_in_2_90),
       .start_out  (start_out_2_90),
       .data_out   (data_out_2_90),
       .op_out     (op_out_2_90),
       .pivot_out  (pivot_out_2_90),
       .r          (r_2_90)
     );

  // row 2, col 91

     reg start_in_2_91;
     wire start_out_2_91;

     reg [1:0] op_in_2_91;
     wire [1:0] op_out_2_91;

     wire r_2_91;

     reg data_in_2_91;
     wire data_out_2_91;

     reg pivot_in_2_91;
     wire pivot_out_2_91;

     always @(posedge clk) begin
         op_in_2_91 <= op_out_2_90;
         pivot_in_2_91 <= pivot_out_2_90;
         start_in_2_91 <= start_out_2_90;
     end

     always @(posedge clk) begin
         data_in_2_91 <= data_out_1_91;
     end
  
     processor_AB AB_2_91 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_91),
       .start_in   (start_in_2_91),
       .op_in      (op_in_2_91),
       .pivot_in   (pivot_in_2_91),
       .start_out  (start_out_2_91),
       .data_out   (data_out_2_91),
       .op_out     (op_out_2_91),
       .pivot_out  (pivot_out_2_91),
       .r          (r_2_91)
     );

  // row 2, col 92

     reg start_in_2_92;
     wire start_out_2_92;

     reg [1:0] op_in_2_92;
     wire [1:0] op_out_2_92;

     wire r_2_92;

     reg data_in_2_92;
     wire data_out_2_92;

     reg pivot_in_2_92;
     wire pivot_out_2_92;

     always @(posedge clk) begin
         op_in_2_92 <= op_out_2_91;
         pivot_in_2_92 <= pivot_out_2_91;
         start_in_2_92 <= start_out_2_91;
     end

     always @(posedge clk) begin
         data_in_2_92 <= data_out_1_92;
     end
  
     processor_AB AB_2_92 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_92),
       .start_in   (start_in_2_92),
       .op_in      (op_in_2_92),
       .pivot_in   (pivot_in_2_92),
       .start_out  (start_out_2_92),
       .data_out   (data_out_2_92),
       .op_out     (op_out_2_92),
       .pivot_out  (pivot_out_2_92),
       .r          (r_2_92)
     );

  // row 2, col 93

     reg start_in_2_93;
     wire start_out_2_93;

     reg [1:0] op_in_2_93;
     wire [1:0] op_out_2_93;

     wire r_2_93;

     reg data_in_2_93;
     wire data_out_2_93;

     reg pivot_in_2_93;
     wire pivot_out_2_93;

     always @(posedge clk) begin
         op_in_2_93 <= op_out_2_92;
         pivot_in_2_93 <= pivot_out_2_92;
         start_in_2_93 <= start_out_2_92;
     end

     always @(posedge clk) begin
         data_in_2_93 <= data_out_1_93;
     end
  
     processor_AB AB_2_93 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_93),
       .start_in   (start_in_2_93),
       .op_in      (op_in_2_93),
       .pivot_in   (pivot_in_2_93),
       .start_out  (start_out_2_93),
       .data_out   (data_out_2_93),
       .op_out     (op_out_2_93),
       .pivot_out  (pivot_out_2_93),
       .r          (r_2_93)
     );

  // row 2, col 94

     reg start_in_2_94;
     wire start_out_2_94;

     reg [1:0] op_in_2_94;
     wire [1:0] op_out_2_94;

     wire r_2_94;

     reg data_in_2_94;
     wire data_out_2_94;

     reg pivot_in_2_94;
     wire pivot_out_2_94;

     always @(posedge clk) begin
         op_in_2_94 <= op_out_2_93;
         pivot_in_2_94 <= pivot_out_2_93;
         start_in_2_94 <= start_out_2_93;
     end

     always @(posedge clk) begin
         data_in_2_94 <= data_out_1_94;
     end
  
     processor_AB AB_2_94 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_94),
       .start_in   (start_in_2_94),
       .op_in      (op_in_2_94),
       .pivot_in   (pivot_in_2_94),
       .start_out  (start_out_2_94),
       .data_out   (data_out_2_94),
       .op_out     (op_out_2_94),
       .pivot_out  (pivot_out_2_94),
       .r          (r_2_94)
     );

  // row 2, col 95

     reg start_in_2_95;
     wire start_out_2_95;

     reg [1:0] op_in_2_95;
     wire [1:0] op_out_2_95;

     wire r_2_95;

     reg data_in_2_95;
     wire data_out_2_95;

     reg pivot_in_2_95;
     wire pivot_out_2_95;

     always @(posedge clk) begin
         op_in_2_95 <= op_out_2_94;
         pivot_in_2_95 <= pivot_out_2_94;
         start_in_2_95 <= start_out_2_94;
     end

     always @(posedge clk) begin
         data_in_2_95 <= data_out_1_95;
     end
  
     processor_AB AB_2_95 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_95),
       .start_in   (start_in_2_95),
       .op_in      (op_in_2_95),
       .pivot_in   (pivot_in_2_95),
       .start_out  (start_out_2_95),
       .data_out   (data_out_2_95),
       .op_out     (op_out_2_95),
       .pivot_out  (pivot_out_2_95),
       .r          (r_2_95)
     );

  // row 2, col 96

     reg start_in_2_96;
     wire start_out_2_96;

     reg [1:0] op_in_2_96;
     wire [1:0] op_out_2_96;

     wire r_2_96;

     reg data_in_2_96;
     wire data_out_2_96;

     reg pivot_in_2_96;
     wire pivot_out_2_96;

     always @(posedge clk) begin
         op_in_2_96 <= op_out_2_95;
         pivot_in_2_96 <= pivot_out_2_95;
         start_in_2_96 <= start_out_2_95;
     end

     always @(posedge clk) begin
         data_in_2_96 <= data_out_1_96;
     end
  
     processor_AB AB_2_96 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_96),
       .start_in   (start_in_2_96),
       .op_in      (op_in_2_96),
       .pivot_in   (pivot_in_2_96),
       .start_out  (start_out_2_96),
       .data_out   (data_out_2_96),
       .op_out     (op_out_2_96),
       .pivot_out  (pivot_out_2_96),
       .r          (r_2_96)
     );

  // row 2, col 97

     reg start_in_2_97;
     wire start_out_2_97;

     reg [1:0] op_in_2_97;
     wire [1:0] op_out_2_97;

     wire r_2_97;

     reg data_in_2_97;
     wire data_out_2_97;

     reg pivot_in_2_97;
     wire pivot_out_2_97;

     always @(posedge clk) begin
         op_in_2_97 <= op_out_2_96;
         pivot_in_2_97 <= pivot_out_2_96;
         start_in_2_97 <= start_out_2_96;
     end

     always @(posedge clk) begin
         data_in_2_97 <= data_out_1_97;
     end
  
     processor_AB AB_2_97 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_97),
       .start_in   (start_in_2_97),
       .op_in      (op_in_2_97),
       .pivot_in   (pivot_in_2_97),
       .start_out  (start_out_2_97),
       .data_out   (data_out_2_97),
       .op_out     (op_out_2_97),
       .pivot_out  (pivot_out_2_97),
       .r          (r_2_97)
     );

  // row 2, col 98

     reg start_in_2_98;
     wire start_out_2_98;

     reg [1:0] op_in_2_98;
     wire [1:0] op_out_2_98;

     wire r_2_98;

     reg data_in_2_98;
     wire data_out_2_98;

     reg pivot_in_2_98;
     wire pivot_out_2_98;

     always @(posedge clk) begin
         op_in_2_98 <= op_out_2_97;
         pivot_in_2_98 <= pivot_out_2_97;
         start_in_2_98 <= start_out_2_97;
     end

     always @(posedge clk) begin
         data_in_2_98 <= data_out_1_98;
     end
  
     processor_AB AB_2_98 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_98),
       .start_in   (start_in_2_98),
       .op_in      (op_in_2_98),
       .pivot_in   (pivot_in_2_98),
       .start_out  (start_out_2_98),
       .data_out   (data_out_2_98),
       .op_out     (op_out_2_98),
       .pivot_out  (pivot_out_2_98),
       .r          (r_2_98)
     );

  // row 2, col 99

     reg start_in_2_99;
     wire start_out_2_99;

     reg [1:0] op_in_2_99;
     wire [1:0] op_out_2_99;

     wire r_2_99;

     reg data_in_2_99;
     wire data_out_2_99;

     reg pivot_in_2_99;
     wire pivot_out_2_99;

     always @(posedge clk) begin
         op_in_2_99 <= op_out_2_98;
         pivot_in_2_99 <= pivot_out_2_98;
         start_in_2_99 <= start_out_2_98;
     end

     always @(posedge clk) begin
         data_in_2_99 <= data_out_1_99;
     end
  
     processor_AB AB_2_99 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_99),
       .start_in   (start_in_2_99),
       .op_in      (op_in_2_99),
       .pivot_in   (pivot_in_2_99),
       .start_out  (start_out_2_99),
       .data_out   (data_out_2_99),
       .op_out     (op_out_2_99),
       .pivot_out  (pivot_out_2_99),
       .r          (r_2_99)
     );

  // row 2, col 100

     reg start_in_2_100;
     wire start_out_2_100;

     reg [1:0] op_in_2_100;
     wire [1:0] op_out_2_100;

     wire r_2_100;

     reg data_in_2_100;
     wire data_out_2_100;

     reg pivot_in_2_100;
     wire pivot_out_2_100;

     always @(posedge clk) begin
         op_in_2_100 <= op_out_2_99;
         pivot_in_2_100 <= pivot_out_2_99;
         start_in_2_100 <= start_out_2_99;
     end

     always @(posedge clk) begin
         data_in_2_100 <= data_out_1_100;
     end
  
     processor_AB AB_2_100 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_100),
       .start_in   (start_in_2_100),
       .op_in      (op_in_2_100),
       .pivot_in   (pivot_in_2_100),
       .start_out  (start_out_2_100),
       .data_out   (data_out_2_100),
       .op_out     (op_out_2_100),
       .pivot_out  (pivot_out_2_100),
       .r          (r_2_100)
     );

  /////////////////////////////////////
  // row 3
  // row 3, col 0

     wire start_in_3_0;
     wire start_out_3_0;

     wire [1:0] op_in_3_0;
     wire [1:0] op_out_3_0;

     wire r_3_0;

     reg data_in_3_0;
     wire data_out_3_0;

     wire pivot_in_3_0;
     wire pivout_out_3_0;

     assign op_in_3_0 = mode & start ? 2'b01 : 2'b00;
     assign pivot_in_3_0 = 0;

     assign start_in_3_0 = start_row[3]; 

     always @(posedge clk) begin
         data_in_3_0 <= data_out_2_0;
     end

     processor_AB AB_3_0 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_0),
       .start_in   (start_in_3_0),
       .op_in      (op_in_3_0),
       .pivot_in   (pivot_in_3_0),
       .start_out  (start_out_3_0),
       .data_out   (data_out_3_0),
       .op_out     (op_out_3_0),
       .pivot_out  (pivot_out_3_0),
       .r          (r_3_0)
     );

  // row 3, col 1

     reg start_in_3_1;
     wire start_out_3_1;

     reg [1:0] op_in_3_1;
     wire [1:0] op_out_3_1;

     wire r_3_1;

     reg data_in_3_1;
     wire data_out_3_1;

     reg pivot_in_3_1;
     wire pivot_out_3_1;

     always @(posedge clk) begin
         op_in_3_1 <= op_out_3_0;
         pivot_in_3_1 <= pivot_out_3_0;
         start_in_3_1 <= start_out_3_0;
     end

     always @(posedge clk) begin
         data_in_3_1 <= data_out_2_1;
     end
  
     processor_AB AB_3_1 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_1),
       .start_in   (start_in_3_1),
       .op_in      (op_in_3_1),
       .pivot_in   (pivot_in_3_1),
       .start_out  (start_out_3_1),
       .data_out   (data_out_3_1),
       .op_out     (op_out_3_1),
       .pivot_out  (pivot_out_3_1),
       .r          (r_3_1)
     );

  // row 3, col 2

     reg start_in_3_2;
     wire start_out_3_2;

     reg [1:0] op_in_3_2;
     wire [1:0] op_out_3_2;

     wire r_3_2;

     reg data_in_3_2;
     wire data_out_3_2;

     reg pivot_in_3_2;
     wire pivot_out_3_2;

     always @(posedge clk) begin
         op_in_3_2 <= op_out_3_1;
         pivot_in_3_2 <= pivot_out_3_1;
         start_in_3_2 <= start_out_3_1;
     end

     always @(posedge clk) begin
         data_in_3_2 <= data_out_2_2;
     end
  
     processor_AB AB_3_2 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_2),
       .start_in   (start_in_3_2),
       .op_in      (op_in_3_2),
       .pivot_in   (pivot_in_3_2),
       .start_out  (start_out_3_2),
       .data_out   (data_out_3_2),
       .op_out     (op_out_3_2),
       .pivot_out  (pivot_out_3_2),
       .r          (r_3_2)
     );

  // row 3, col 3

     reg start_in_3_3;
     wire start_out_3_3;

     reg [1:0] op_in_3_3;
     wire [1:0] op_out_3_3;

     wire r_3_3;

     reg data_in_3_3;
     wire data_out_3_3;

     reg pivot_in_3_3;
     wire pivot_out_3_3;

     always @(posedge clk) begin
         op_in_3_3 <= op_out_3_2;
         pivot_in_3_3 <= pivot_out_3_2;
         start_in_3_3 <= start_out_3_2;
     end

     always @(posedge clk) begin
         data_in_3_3 <= data_out_2_3;
     end
  
     processor_AB AB_3_3 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_3),
       .start_in   (start_in_3_3),
       .op_in      (op_in_3_3),
       .pivot_in   (pivot_in_3_3),
       .start_out  (start_out_3_3),
       .data_out   (data_out_3_3),
       .op_out     (op_out_3_3),
       .pivot_out  (pivot_out_3_3),
       .r          (r_3_3)
     );

  // row 3, col 4

     reg start_in_3_4;
     wire start_out_3_4;

     reg [1:0] op_in_3_4;
     wire [1:0] op_out_3_4;

     wire r_3_4;

     reg data_in_3_4;
     wire data_out_3_4;

     reg pivot_in_3_4;
     wire pivot_out_3_4;

     always @(posedge clk) begin
         op_in_3_4 <= op_out_3_3;
         pivot_in_3_4 <= pivot_out_3_3;
         start_in_3_4 <= start_out_3_3;
     end

     always @(posedge clk) begin
         data_in_3_4 <= data_out_2_4;
     end
  
     processor_AB AB_3_4 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_4),
       .start_in   (start_in_3_4),
       .op_in      (op_in_3_4),
       .pivot_in   (pivot_in_3_4),
       .start_out  (start_out_3_4),
       .data_out   (data_out_3_4),
       .op_out     (op_out_3_4),
       .pivot_out  (pivot_out_3_4),
       .r          (r_3_4)
     );

  // row 3, col 5

     reg start_in_3_5;
     wire start_out_3_5;

     reg [1:0] op_in_3_5;
     wire [1:0] op_out_3_5;

     wire r_3_5;

     reg data_in_3_5;
     wire data_out_3_5;

     reg pivot_in_3_5;
     wire pivot_out_3_5;

     always @(posedge clk) begin
         op_in_3_5 <= op_out_3_4;
         pivot_in_3_5 <= pivot_out_3_4;
         start_in_3_5 <= start_out_3_4;
     end

     always @(posedge clk) begin
         data_in_3_5 <= data_out_2_5;
     end
  
     processor_AB AB_3_5 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_5),
       .start_in   (start_in_3_5),
       .op_in      (op_in_3_5),
       .pivot_in   (pivot_in_3_5),
       .start_out  (start_out_3_5),
       .data_out   (data_out_3_5),
       .op_out     (op_out_3_5),
       .pivot_out  (pivot_out_3_5),
       .r          (r_3_5)
     );

  // row 3, col 6

     reg start_in_3_6;
     wire start_out_3_6;

     reg [1:0] op_in_3_6;
     wire [1:0] op_out_3_6;

     wire r_3_6;

     reg data_in_3_6;
     wire data_out_3_6;

     reg pivot_in_3_6;
     wire pivot_out_3_6;

     always @(posedge clk) begin
         op_in_3_6 <= op_out_3_5;
         pivot_in_3_6 <= pivot_out_3_5;
         start_in_3_6 <= start_out_3_5;
     end

     always @(posedge clk) begin
         data_in_3_6 <= data_out_2_6;
     end
  
     processor_AB AB_3_6 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_6),
       .start_in   (start_in_3_6),
       .op_in      (op_in_3_6),
       .pivot_in   (pivot_in_3_6),
       .start_out  (start_out_3_6),
       .data_out   (data_out_3_6),
       .op_out     (op_out_3_6),
       .pivot_out  (pivot_out_3_6),
       .r          (r_3_6)
     );

  // row 3, col 7

     reg start_in_3_7;
     wire start_out_3_7;

     reg [1:0] op_in_3_7;
     wire [1:0] op_out_3_7;

     wire r_3_7;

     reg data_in_3_7;
     wire data_out_3_7;

     reg pivot_in_3_7;
     wire pivot_out_3_7;

     always @(posedge clk) begin
         op_in_3_7 <= op_out_3_6;
         pivot_in_3_7 <= pivot_out_3_6;
         start_in_3_7 <= start_out_3_6;
     end

     always @(posedge clk) begin
         data_in_3_7 <= data_out_2_7;
     end
  
     processor_AB AB_3_7 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_7),
       .start_in   (start_in_3_7),
       .op_in      (op_in_3_7),
       .pivot_in   (pivot_in_3_7),
       .start_out  (start_out_3_7),
       .data_out   (data_out_3_7),
       .op_out     (op_out_3_7),
       .pivot_out  (pivot_out_3_7),
       .r          (r_3_7)
     );

  // row 3, col 8

     reg start_in_3_8;
     wire start_out_3_8;

     reg [1:0] op_in_3_8;
     wire [1:0] op_out_3_8;

     wire r_3_8;

     reg data_in_3_8;
     wire data_out_3_8;

     reg pivot_in_3_8;
     wire pivot_out_3_8;

     always @(posedge clk) begin
         op_in_3_8 <= op_out_3_7;
         pivot_in_3_8 <= pivot_out_3_7;
         start_in_3_8 <= start_out_3_7;
     end

     always @(posedge clk) begin
         data_in_3_8 <= data_out_2_8;
     end
  
     processor_AB AB_3_8 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_8),
       .start_in   (start_in_3_8),
       .op_in      (op_in_3_8),
       .pivot_in   (pivot_in_3_8),
       .start_out  (start_out_3_8),
       .data_out   (data_out_3_8),
       .op_out     (op_out_3_8),
       .pivot_out  (pivot_out_3_8),
       .r          (r_3_8)
     );

  // row 3, col 9

     reg start_in_3_9;
     wire start_out_3_9;

     reg [1:0] op_in_3_9;
     wire [1:0] op_out_3_9;

     wire r_3_9;

     reg data_in_3_9;
     wire data_out_3_9;

     reg pivot_in_3_9;
     wire pivot_out_3_9;

     always @(posedge clk) begin
         op_in_3_9 <= op_out_3_8;
         pivot_in_3_9 <= pivot_out_3_8;
         start_in_3_9 <= start_out_3_8;
     end

     always @(posedge clk) begin
         data_in_3_9 <= data_out_2_9;
     end
  
     processor_AB AB_3_9 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_9),
       .start_in   (start_in_3_9),
       .op_in      (op_in_3_9),
       .pivot_in   (pivot_in_3_9),
       .start_out  (start_out_3_9),
       .data_out   (data_out_3_9),
       .op_out     (op_out_3_9),
       .pivot_out  (pivot_out_3_9),
       .r          (r_3_9)
     );

  // row 3, col 10

     reg start_in_3_10;
     wire start_out_3_10;

     reg [1:0] op_in_3_10;
     wire [1:0] op_out_3_10;

     wire r_3_10;

     reg data_in_3_10;
     wire data_out_3_10;

     reg pivot_in_3_10;
     wire pivot_out_3_10;

     always @(posedge clk) begin
         op_in_3_10 <= op_out_3_9;
         pivot_in_3_10 <= pivot_out_3_9;
         start_in_3_10 <= start_out_3_9;
     end

     always @(posedge clk) begin
         data_in_3_10 <= data_out_2_10;
     end
  
     processor_AB AB_3_10 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_10),
       .start_in   (start_in_3_10),
       .op_in      (op_in_3_10),
       .pivot_in   (pivot_in_3_10),
       .start_out  (start_out_3_10),
       .data_out   (data_out_3_10),
       .op_out     (op_out_3_10),
       .pivot_out  (pivot_out_3_10),
       .r          (r_3_10)
     );

  // row 3, col 11

     reg start_in_3_11;
     wire start_out_3_11;

     reg [1:0] op_in_3_11;
     wire [1:0] op_out_3_11;

     wire r_3_11;

     reg data_in_3_11;
     wire data_out_3_11;

     reg pivot_in_3_11;
     wire pivot_out_3_11;

     always @(posedge clk) begin
         op_in_3_11 <= op_out_3_10;
         pivot_in_3_11 <= pivot_out_3_10;
         start_in_3_11 <= start_out_3_10;
     end

     always @(posedge clk) begin
         data_in_3_11 <= data_out_2_11;
     end
  
     processor_AB AB_3_11 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_11),
       .start_in   (start_in_3_11),
       .op_in      (op_in_3_11),
       .pivot_in   (pivot_in_3_11),
       .start_out  (start_out_3_11),
       .data_out   (data_out_3_11),
       .op_out     (op_out_3_11),
       .pivot_out  (pivot_out_3_11),
       .r          (r_3_11)
     );

  // row 3, col 12

     reg start_in_3_12;
     wire start_out_3_12;

     reg [1:0] op_in_3_12;
     wire [1:0] op_out_3_12;

     wire r_3_12;

     reg data_in_3_12;
     wire data_out_3_12;

     reg pivot_in_3_12;
     wire pivot_out_3_12;

     always @(posedge clk) begin
         op_in_3_12 <= op_out_3_11;
         pivot_in_3_12 <= pivot_out_3_11;
         start_in_3_12 <= start_out_3_11;
     end

     always @(posedge clk) begin
         data_in_3_12 <= data_out_2_12;
     end
  
     processor_AB AB_3_12 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_12),
       .start_in   (start_in_3_12),
       .op_in      (op_in_3_12),
       .pivot_in   (pivot_in_3_12),
       .start_out  (start_out_3_12),
       .data_out   (data_out_3_12),
       .op_out     (op_out_3_12),
       .pivot_out  (pivot_out_3_12),
       .r          (r_3_12)
     );

  // row 3, col 13

     reg start_in_3_13;
     wire start_out_3_13;

     reg [1:0] op_in_3_13;
     wire [1:0] op_out_3_13;

     wire r_3_13;

     reg data_in_3_13;
     wire data_out_3_13;

     reg pivot_in_3_13;
     wire pivot_out_3_13;

     always @(posedge clk) begin
         op_in_3_13 <= op_out_3_12;
         pivot_in_3_13 <= pivot_out_3_12;
         start_in_3_13 <= start_out_3_12;
     end

     always @(posedge clk) begin
         data_in_3_13 <= data_out_2_13;
     end
  
     processor_AB AB_3_13 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_13),
       .start_in   (start_in_3_13),
       .op_in      (op_in_3_13),
       .pivot_in   (pivot_in_3_13),
       .start_out  (start_out_3_13),
       .data_out   (data_out_3_13),
       .op_out     (op_out_3_13),
       .pivot_out  (pivot_out_3_13),
       .r          (r_3_13)
     );

  // row 3, col 14

     reg start_in_3_14;
     wire start_out_3_14;

     reg [1:0] op_in_3_14;
     wire [1:0] op_out_3_14;

     wire r_3_14;

     reg data_in_3_14;
     wire data_out_3_14;

     reg pivot_in_3_14;
     wire pivot_out_3_14;

     always @(posedge clk) begin
         op_in_3_14 <= op_out_3_13;
         pivot_in_3_14 <= pivot_out_3_13;
         start_in_3_14 <= start_out_3_13;
     end

     always @(posedge clk) begin
         data_in_3_14 <= data_out_2_14;
     end
  
     processor_AB AB_3_14 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_14),
       .start_in   (start_in_3_14),
       .op_in      (op_in_3_14),
       .pivot_in   (pivot_in_3_14),
       .start_out  (start_out_3_14),
       .data_out   (data_out_3_14),
       .op_out     (op_out_3_14),
       .pivot_out  (pivot_out_3_14),
       .r          (r_3_14)
     );

  // row 3, col 15

     reg start_in_3_15;
     wire start_out_3_15;

     reg [1:0] op_in_3_15;
     wire [1:0] op_out_3_15;

     wire r_3_15;

     reg data_in_3_15;
     wire data_out_3_15;

     reg pivot_in_3_15;
     wire pivot_out_3_15;

     always @(posedge clk) begin
         op_in_3_15 <= op_out_3_14;
         pivot_in_3_15 <= pivot_out_3_14;
         start_in_3_15 <= start_out_3_14;
     end

     always @(posedge clk) begin
         data_in_3_15 <= data_out_2_15;
     end
  
     processor_AB AB_3_15 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_15),
       .start_in   (start_in_3_15),
       .op_in      (op_in_3_15),
       .pivot_in   (pivot_in_3_15),
       .start_out  (start_out_3_15),
       .data_out   (data_out_3_15),
       .op_out     (op_out_3_15),
       .pivot_out  (pivot_out_3_15),
       .r          (r_3_15)
     );

  // row 3, col 16

     reg start_in_3_16;
     wire start_out_3_16;

     reg [1:0] op_in_3_16;
     wire [1:0] op_out_3_16;

     wire r_3_16;

     reg data_in_3_16;
     wire data_out_3_16;

     reg pivot_in_3_16;
     wire pivot_out_3_16;

     always @(posedge clk) begin
         op_in_3_16 <= op_out_3_15;
         pivot_in_3_16 <= pivot_out_3_15;
         start_in_3_16 <= start_out_3_15;
     end

     always @(posedge clk) begin
         data_in_3_16 <= data_out_2_16;
     end
  
     processor_AB AB_3_16 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_16),
       .start_in   (start_in_3_16),
       .op_in      (op_in_3_16),
       .pivot_in   (pivot_in_3_16),
       .start_out  (start_out_3_16),
       .data_out   (data_out_3_16),
       .op_out     (op_out_3_16),
       .pivot_out  (pivot_out_3_16),
       .r          (r_3_16)
     );

  // row 3, col 17

     reg start_in_3_17;
     wire start_out_3_17;

     reg [1:0] op_in_3_17;
     wire [1:0] op_out_3_17;

     wire r_3_17;

     reg data_in_3_17;
     wire data_out_3_17;

     reg pivot_in_3_17;
     wire pivot_out_3_17;

     always @(posedge clk) begin
         op_in_3_17 <= op_out_3_16;
         pivot_in_3_17 <= pivot_out_3_16;
         start_in_3_17 <= start_out_3_16;
     end

     always @(posedge clk) begin
         data_in_3_17 <= data_out_2_17;
     end
  
     processor_AB AB_3_17 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_17),
       .start_in   (start_in_3_17),
       .op_in      (op_in_3_17),
       .pivot_in   (pivot_in_3_17),
       .start_out  (start_out_3_17),
       .data_out   (data_out_3_17),
       .op_out     (op_out_3_17),
       .pivot_out  (pivot_out_3_17),
       .r          (r_3_17)
     );

  // row 3, col 18

     reg start_in_3_18;
     wire start_out_3_18;

     reg [1:0] op_in_3_18;
     wire [1:0] op_out_3_18;

     wire r_3_18;

     reg data_in_3_18;
     wire data_out_3_18;

     reg pivot_in_3_18;
     wire pivot_out_3_18;

     always @(posedge clk) begin
         op_in_3_18 <= op_out_3_17;
         pivot_in_3_18 <= pivot_out_3_17;
         start_in_3_18 <= start_out_3_17;
     end

     always @(posedge clk) begin
         data_in_3_18 <= data_out_2_18;
     end
  
     processor_AB AB_3_18 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_18),
       .start_in   (start_in_3_18),
       .op_in      (op_in_3_18),
       .pivot_in   (pivot_in_3_18),
       .start_out  (start_out_3_18),
       .data_out   (data_out_3_18),
       .op_out     (op_out_3_18),
       .pivot_out  (pivot_out_3_18),
       .r          (r_3_18)
     );

  // row 3, col 19

     reg start_in_3_19;
     wire start_out_3_19;

     reg [1:0] op_in_3_19;
     wire [1:0] op_out_3_19;

     wire r_3_19;

     reg data_in_3_19;
     wire data_out_3_19;

     reg pivot_in_3_19;
     wire pivot_out_3_19;

     always @(posedge clk) begin
         op_in_3_19 <= op_out_3_18;
         pivot_in_3_19 <= pivot_out_3_18;
         start_in_3_19 <= start_out_3_18;
     end

     always @(posedge clk) begin
         data_in_3_19 <= data_out_2_19;
     end
  
     processor_AB AB_3_19 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_19),
       .start_in   (start_in_3_19),
       .op_in      (op_in_3_19),
       .pivot_in   (pivot_in_3_19),
       .start_out  (start_out_3_19),
       .data_out   (data_out_3_19),
       .op_out     (op_out_3_19),
       .pivot_out  (pivot_out_3_19),
       .r          (r_3_19)
     );

  // row 3, col 20

     reg start_in_3_20;
     wire start_out_3_20;

     reg [1:0] op_in_3_20;
     wire [1:0] op_out_3_20;

     wire r_3_20;

     reg data_in_3_20;
     wire data_out_3_20;

     reg pivot_in_3_20;
     wire pivot_out_3_20;

     always @(posedge clk) begin
         op_in_3_20 <= op_out_3_19;
         pivot_in_3_20 <= pivot_out_3_19;
         start_in_3_20 <= start_out_3_19;
     end

     always @(posedge clk) begin
         data_in_3_20 <= data_out_2_20;
     end
  
     processor_AB AB_3_20 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_20),
       .start_in   (start_in_3_20),
       .op_in      (op_in_3_20),
       .pivot_in   (pivot_in_3_20),
       .start_out  (start_out_3_20),
       .data_out   (data_out_3_20),
       .op_out     (op_out_3_20),
       .pivot_out  (pivot_out_3_20),
       .r          (r_3_20)
     );

  // row 3, col 21

     reg start_in_3_21;
     wire start_out_3_21;

     reg [1:0] op_in_3_21;
     wire [1:0] op_out_3_21;

     wire r_3_21;

     reg data_in_3_21;
     wire data_out_3_21;

     reg pivot_in_3_21;
     wire pivot_out_3_21;

     always @(posedge clk) begin
         op_in_3_21 <= op_out_3_20;
         pivot_in_3_21 <= pivot_out_3_20;
         start_in_3_21 <= start_out_3_20;
     end

     always @(posedge clk) begin
         data_in_3_21 <= data_out_2_21;
     end
  
     processor_AB AB_3_21 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_21),
       .start_in   (start_in_3_21),
       .op_in      (op_in_3_21),
       .pivot_in   (pivot_in_3_21),
       .start_out  (start_out_3_21),
       .data_out   (data_out_3_21),
       .op_out     (op_out_3_21),
       .pivot_out  (pivot_out_3_21),
       .r          (r_3_21)
     );

  // row 3, col 22

     reg start_in_3_22;
     wire start_out_3_22;

     reg [1:0] op_in_3_22;
     wire [1:0] op_out_3_22;

     wire r_3_22;

     reg data_in_3_22;
     wire data_out_3_22;

     reg pivot_in_3_22;
     wire pivot_out_3_22;

     always @(posedge clk) begin
         op_in_3_22 <= op_out_3_21;
         pivot_in_3_22 <= pivot_out_3_21;
         start_in_3_22 <= start_out_3_21;
     end

     always @(posedge clk) begin
         data_in_3_22 <= data_out_2_22;
     end
  
     processor_AB AB_3_22 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_22),
       .start_in   (start_in_3_22),
       .op_in      (op_in_3_22),
       .pivot_in   (pivot_in_3_22),
       .start_out  (start_out_3_22),
       .data_out   (data_out_3_22),
       .op_out     (op_out_3_22),
       .pivot_out  (pivot_out_3_22),
       .r          (r_3_22)
     );

  // row 3, col 23

     reg start_in_3_23;
     wire start_out_3_23;

     reg [1:0] op_in_3_23;
     wire [1:0] op_out_3_23;

     wire r_3_23;

     reg data_in_3_23;
     wire data_out_3_23;

     reg pivot_in_3_23;
     wire pivot_out_3_23;

     always @(posedge clk) begin
         op_in_3_23 <= op_out_3_22;
         pivot_in_3_23 <= pivot_out_3_22;
         start_in_3_23 <= start_out_3_22;
     end

     always @(posedge clk) begin
         data_in_3_23 <= data_out_2_23;
     end
  
     processor_AB AB_3_23 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_23),
       .start_in   (start_in_3_23),
       .op_in      (op_in_3_23),
       .pivot_in   (pivot_in_3_23),
       .start_out  (start_out_3_23),
       .data_out   (data_out_3_23),
       .op_out     (op_out_3_23),
       .pivot_out  (pivot_out_3_23),
       .r          (r_3_23)
     );

  // row 3, col 24

     reg start_in_3_24;
     wire start_out_3_24;

     reg [1:0] op_in_3_24;
     wire [1:0] op_out_3_24;

     wire r_3_24;

     reg data_in_3_24;
     wire data_out_3_24;

     reg pivot_in_3_24;
     wire pivot_out_3_24;

     always @(posedge clk) begin
         op_in_3_24 <= op_out_3_23;
         pivot_in_3_24 <= pivot_out_3_23;
         start_in_3_24 <= start_out_3_23;
     end

     always @(posedge clk) begin
         data_in_3_24 <= data_out_2_24;
     end
  
     processor_AB AB_3_24 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_24),
       .start_in   (start_in_3_24),
       .op_in      (op_in_3_24),
       .pivot_in   (pivot_in_3_24),
       .start_out  (start_out_3_24),
       .data_out   (data_out_3_24),
       .op_out     (op_out_3_24),
       .pivot_out  (pivot_out_3_24),
       .r          (r_3_24)
     );

  // row 3, col 25

     reg start_in_3_25;
     wire start_out_3_25;

     reg [1:0] op_in_3_25;
     wire [1:0] op_out_3_25;

     wire r_3_25;

     reg data_in_3_25;
     wire data_out_3_25;

     reg pivot_in_3_25;
     wire pivot_out_3_25;

     always @(posedge clk) begin
         op_in_3_25 <= op_out_3_24;
         pivot_in_3_25 <= pivot_out_3_24;
         start_in_3_25 <= start_out_3_24;
     end

     always @(posedge clk) begin
         data_in_3_25 <= data_out_2_25;
     end
  
     processor_AB AB_3_25 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_25),
       .start_in   (start_in_3_25),
       .op_in      (op_in_3_25),
       .pivot_in   (pivot_in_3_25),
       .start_out  (start_out_3_25),
       .data_out   (data_out_3_25),
       .op_out     (op_out_3_25),
       .pivot_out  (pivot_out_3_25),
       .r          (r_3_25)
     );

  // row 3, col 26

     reg start_in_3_26;
     wire start_out_3_26;

     reg [1:0] op_in_3_26;
     wire [1:0] op_out_3_26;

     wire r_3_26;

     reg data_in_3_26;
     wire data_out_3_26;

     reg pivot_in_3_26;
     wire pivot_out_3_26;

     always @(posedge clk) begin
         op_in_3_26 <= op_out_3_25;
         pivot_in_3_26 <= pivot_out_3_25;
         start_in_3_26 <= start_out_3_25;
     end

     always @(posedge clk) begin
         data_in_3_26 <= data_out_2_26;
     end
  
     processor_AB AB_3_26 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_26),
       .start_in   (start_in_3_26),
       .op_in      (op_in_3_26),
       .pivot_in   (pivot_in_3_26),
       .start_out  (start_out_3_26),
       .data_out   (data_out_3_26),
       .op_out     (op_out_3_26),
       .pivot_out  (pivot_out_3_26),
       .r          (r_3_26)
     );

  // row 3, col 27

     reg start_in_3_27;
     wire start_out_3_27;

     reg [1:0] op_in_3_27;
     wire [1:0] op_out_3_27;

     wire r_3_27;

     reg data_in_3_27;
     wire data_out_3_27;

     reg pivot_in_3_27;
     wire pivot_out_3_27;

     always @(posedge clk) begin
         op_in_3_27 <= op_out_3_26;
         pivot_in_3_27 <= pivot_out_3_26;
         start_in_3_27 <= start_out_3_26;
     end

     always @(posedge clk) begin
         data_in_3_27 <= data_out_2_27;
     end
  
     processor_AB AB_3_27 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_27),
       .start_in   (start_in_3_27),
       .op_in      (op_in_3_27),
       .pivot_in   (pivot_in_3_27),
       .start_out  (start_out_3_27),
       .data_out   (data_out_3_27),
       .op_out     (op_out_3_27),
       .pivot_out  (pivot_out_3_27),
       .r          (r_3_27)
     );

  // row 3, col 28

     reg start_in_3_28;
     wire start_out_3_28;

     reg [1:0] op_in_3_28;
     wire [1:0] op_out_3_28;

     wire r_3_28;

     reg data_in_3_28;
     wire data_out_3_28;

     reg pivot_in_3_28;
     wire pivot_out_3_28;

     always @(posedge clk) begin
         op_in_3_28 <= op_out_3_27;
         pivot_in_3_28 <= pivot_out_3_27;
         start_in_3_28 <= start_out_3_27;
     end

     always @(posedge clk) begin
         data_in_3_28 <= data_out_2_28;
     end
  
     processor_AB AB_3_28 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_28),
       .start_in   (start_in_3_28),
       .op_in      (op_in_3_28),
       .pivot_in   (pivot_in_3_28),
       .start_out  (start_out_3_28),
       .data_out   (data_out_3_28),
       .op_out     (op_out_3_28),
       .pivot_out  (pivot_out_3_28),
       .r          (r_3_28)
     );

  // row 3, col 29

     reg start_in_3_29;
     wire start_out_3_29;

     reg [1:0] op_in_3_29;
     wire [1:0] op_out_3_29;

     wire r_3_29;

     reg data_in_3_29;
     wire data_out_3_29;

     reg pivot_in_3_29;
     wire pivot_out_3_29;

     always @(posedge clk) begin
         op_in_3_29 <= op_out_3_28;
         pivot_in_3_29 <= pivot_out_3_28;
         start_in_3_29 <= start_out_3_28;
     end

     always @(posedge clk) begin
         data_in_3_29 <= data_out_2_29;
     end
  
     processor_AB AB_3_29 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_29),
       .start_in   (start_in_3_29),
       .op_in      (op_in_3_29),
       .pivot_in   (pivot_in_3_29),
       .start_out  (start_out_3_29),
       .data_out   (data_out_3_29),
       .op_out     (op_out_3_29),
       .pivot_out  (pivot_out_3_29),
       .r          (r_3_29)
     );

  // row 3, col 30

     reg start_in_3_30;
     wire start_out_3_30;

     reg [1:0] op_in_3_30;
     wire [1:0] op_out_3_30;

     wire r_3_30;

     reg data_in_3_30;
     wire data_out_3_30;

     reg pivot_in_3_30;
     wire pivot_out_3_30;

     always @(posedge clk) begin
         op_in_3_30 <= op_out_3_29;
         pivot_in_3_30 <= pivot_out_3_29;
         start_in_3_30 <= start_out_3_29;
     end

     always @(posedge clk) begin
         data_in_3_30 <= data_out_2_30;
     end
  
     processor_AB AB_3_30 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_30),
       .start_in   (start_in_3_30),
       .op_in      (op_in_3_30),
       .pivot_in   (pivot_in_3_30),
       .start_out  (start_out_3_30),
       .data_out   (data_out_3_30),
       .op_out     (op_out_3_30),
       .pivot_out  (pivot_out_3_30),
       .r          (r_3_30)
     );

  // row 3, col 31

     reg start_in_3_31;
     wire start_out_3_31;

     reg [1:0] op_in_3_31;
     wire [1:0] op_out_3_31;

     wire r_3_31;

     reg data_in_3_31;
     wire data_out_3_31;

     reg pivot_in_3_31;
     wire pivot_out_3_31;

     always @(posedge clk) begin
         op_in_3_31 <= op_out_3_30;
         pivot_in_3_31 <= pivot_out_3_30;
         start_in_3_31 <= start_out_3_30;
     end

     always @(posedge clk) begin
         data_in_3_31 <= data_out_2_31;
     end
  
     processor_AB AB_3_31 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_31),
       .start_in   (start_in_3_31),
       .op_in      (op_in_3_31),
       .pivot_in   (pivot_in_3_31),
       .start_out  (start_out_3_31),
       .data_out   (data_out_3_31),
       .op_out     (op_out_3_31),
       .pivot_out  (pivot_out_3_31),
       .r          (r_3_31)
     );

  // row 3, col 32

     reg start_in_3_32;
     wire start_out_3_32;

     reg [1:0] op_in_3_32;
     wire [1:0] op_out_3_32;

     wire r_3_32;

     reg data_in_3_32;
     wire data_out_3_32;

     reg pivot_in_3_32;
     wire pivot_out_3_32;

     always @(posedge clk) begin
         op_in_3_32 <= op_out_3_31;
         pivot_in_3_32 <= pivot_out_3_31;
         start_in_3_32 <= start_out_3_31;
     end

     always @(posedge clk) begin
         data_in_3_32 <= data_out_2_32;
     end
  
     processor_AB AB_3_32 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_32),
       .start_in   (start_in_3_32),
       .op_in      (op_in_3_32),
       .pivot_in   (pivot_in_3_32),
       .start_out  (start_out_3_32),
       .data_out   (data_out_3_32),
       .op_out     (op_out_3_32),
       .pivot_out  (pivot_out_3_32),
       .r          (r_3_32)
     );

  // row 3, col 33

     reg start_in_3_33;
     wire start_out_3_33;

     reg [1:0] op_in_3_33;
     wire [1:0] op_out_3_33;

     wire r_3_33;

     reg data_in_3_33;
     wire data_out_3_33;

     reg pivot_in_3_33;
     wire pivot_out_3_33;

     always @(posedge clk) begin
         op_in_3_33 <= op_out_3_32;
         pivot_in_3_33 <= pivot_out_3_32;
         start_in_3_33 <= start_out_3_32;
     end

     always @(posedge clk) begin
         data_in_3_33 <= data_out_2_33;
     end
  
     processor_AB AB_3_33 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_33),
       .start_in   (start_in_3_33),
       .op_in      (op_in_3_33),
       .pivot_in   (pivot_in_3_33),
       .start_out  (start_out_3_33),
       .data_out   (data_out_3_33),
       .op_out     (op_out_3_33),
       .pivot_out  (pivot_out_3_33),
       .r          (r_3_33)
     );

  // row 3, col 34

     reg start_in_3_34;
     wire start_out_3_34;

     reg [1:0] op_in_3_34;
     wire [1:0] op_out_3_34;

     wire r_3_34;

     reg data_in_3_34;
     wire data_out_3_34;

     reg pivot_in_3_34;
     wire pivot_out_3_34;

     always @(posedge clk) begin
         op_in_3_34 <= op_out_3_33;
         pivot_in_3_34 <= pivot_out_3_33;
         start_in_3_34 <= start_out_3_33;
     end

     always @(posedge clk) begin
         data_in_3_34 <= data_out_2_34;
     end
  
     processor_AB AB_3_34 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_34),
       .start_in   (start_in_3_34),
       .op_in      (op_in_3_34),
       .pivot_in   (pivot_in_3_34),
       .start_out  (start_out_3_34),
       .data_out   (data_out_3_34),
       .op_out     (op_out_3_34),
       .pivot_out  (pivot_out_3_34),
       .r          (r_3_34)
     );

  // row 3, col 35

     reg start_in_3_35;
     wire start_out_3_35;

     reg [1:0] op_in_3_35;
     wire [1:0] op_out_3_35;

     wire r_3_35;

     reg data_in_3_35;
     wire data_out_3_35;

     reg pivot_in_3_35;
     wire pivot_out_3_35;

     always @(posedge clk) begin
         op_in_3_35 <= op_out_3_34;
         pivot_in_3_35 <= pivot_out_3_34;
         start_in_3_35 <= start_out_3_34;
     end

     always @(posedge clk) begin
         data_in_3_35 <= data_out_2_35;
     end
  
     processor_AB AB_3_35 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_35),
       .start_in   (start_in_3_35),
       .op_in      (op_in_3_35),
       .pivot_in   (pivot_in_3_35),
       .start_out  (start_out_3_35),
       .data_out   (data_out_3_35),
       .op_out     (op_out_3_35),
       .pivot_out  (pivot_out_3_35),
       .r          (r_3_35)
     );

  // row 3, col 36

     reg start_in_3_36;
     wire start_out_3_36;

     reg [1:0] op_in_3_36;
     wire [1:0] op_out_3_36;

     wire r_3_36;

     reg data_in_3_36;
     wire data_out_3_36;

     reg pivot_in_3_36;
     wire pivot_out_3_36;

     always @(posedge clk) begin
         op_in_3_36 <= op_out_3_35;
         pivot_in_3_36 <= pivot_out_3_35;
         start_in_3_36 <= start_out_3_35;
     end

     always @(posedge clk) begin
         data_in_3_36 <= data_out_2_36;
     end
  
     processor_AB AB_3_36 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_36),
       .start_in   (start_in_3_36),
       .op_in      (op_in_3_36),
       .pivot_in   (pivot_in_3_36),
       .start_out  (start_out_3_36),
       .data_out   (data_out_3_36),
       .op_out     (op_out_3_36),
       .pivot_out  (pivot_out_3_36),
       .r          (r_3_36)
     );

  // row 3, col 37

     reg start_in_3_37;
     wire start_out_3_37;

     reg [1:0] op_in_3_37;
     wire [1:0] op_out_3_37;

     wire r_3_37;

     reg data_in_3_37;
     wire data_out_3_37;

     reg pivot_in_3_37;
     wire pivot_out_3_37;

     always @(posedge clk) begin
         op_in_3_37 <= op_out_3_36;
         pivot_in_3_37 <= pivot_out_3_36;
         start_in_3_37 <= start_out_3_36;
     end

     always @(posedge clk) begin
         data_in_3_37 <= data_out_2_37;
     end
  
     processor_AB AB_3_37 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_37),
       .start_in   (start_in_3_37),
       .op_in      (op_in_3_37),
       .pivot_in   (pivot_in_3_37),
       .start_out  (start_out_3_37),
       .data_out   (data_out_3_37),
       .op_out     (op_out_3_37),
       .pivot_out  (pivot_out_3_37),
       .r          (r_3_37)
     );

  // row 3, col 38

     reg start_in_3_38;
     wire start_out_3_38;

     reg [1:0] op_in_3_38;
     wire [1:0] op_out_3_38;

     wire r_3_38;

     reg data_in_3_38;
     wire data_out_3_38;

     reg pivot_in_3_38;
     wire pivot_out_3_38;

     always @(posedge clk) begin
         op_in_3_38 <= op_out_3_37;
         pivot_in_3_38 <= pivot_out_3_37;
         start_in_3_38 <= start_out_3_37;
     end

     always @(posedge clk) begin
         data_in_3_38 <= data_out_2_38;
     end
  
     processor_AB AB_3_38 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_38),
       .start_in   (start_in_3_38),
       .op_in      (op_in_3_38),
       .pivot_in   (pivot_in_3_38),
       .start_out  (start_out_3_38),
       .data_out   (data_out_3_38),
       .op_out     (op_out_3_38),
       .pivot_out  (pivot_out_3_38),
       .r          (r_3_38)
     );

  // row 3, col 39

     reg start_in_3_39;
     wire start_out_3_39;

     reg [1:0] op_in_3_39;
     wire [1:0] op_out_3_39;

     wire r_3_39;

     reg data_in_3_39;
     wire data_out_3_39;

     reg pivot_in_3_39;
     wire pivot_out_3_39;

     always @(posedge clk) begin
         op_in_3_39 <= op_out_3_38;
         pivot_in_3_39 <= pivot_out_3_38;
         start_in_3_39 <= start_out_3_38;
     end

     always @(posedge clk) begin
         data_in_3_39 <= data_out_2_39;
     end
  
     processor_AB AB_3_39 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_39),
       .start_in   (start_in_3_39),
       .op_in      (op_in_3_39),
       .pivot_in   (pivot_in_3_39),
       .start_out  (start_out_3_39),
       .data_out   (data_out_3_39),
       .op_out     (op_out_3_39),
       .pivot_out  (pivot_out_3_39),
       .r          (r_3_39)
     );

  // row 3, col 40

     reg start_in_3_40;
     wire start_out_3_40;

     reg [1:0] op_in_3_40;
     wire [1:0] op_out_3_40;

     wire r_3_40;

     reg data_in_3_40;
     wire data_out_3_40;

     reg pivot_in_3_40;
     wire pivot_out_3_40;

     always @(posedge clk) begin
         op_in_3_40 <= op_out_3_39;
         pivot_in_3_40 <= pivot_out_3_39;
         start_in_3_40 <= start_out_3_39;
     end

     always @(posedge clk) begin
         data_in_3_40 <= data_out_2_40;
     end
  
     processor_AB AB_3_40 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_40),
       .start_in   (start_in_3_40),
       .op_in      (op_in_3_40),
       .pivot_in   (pivot_in_3_40),
       .start_out  (start_out_3_40),
       .data_out   (data_out_3_40),
       .op_out     (op_out_3_40),
       .pivot_out  (pivot_out_3_40),
       .r          (r_3_40)
     );

  // row 3, col 41

     reg start_in_3_41;
     wire start_out_3_41;

     reg [1:0] op_in_3_41;
     wire [1:0] op_out_3_41;

     wire r_3_41;

     reg data_in_3_41;
     wire data_out_3_41;

     reg pivot_in_3_41;
     wire pivot_out_3_41;

     always @(posedge clk) begin
         op_in_3_41 <= op_out_3_40;
         pivot_in_3_41 <= pivot_out_3_40;
         start_in_3_41 <= start_out_3_40;
     end

     always @(posedge clk) begin
         data_in_3_41 <= data_out_2_41;
     end
  
     processor_AB AB_3_41 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_41),
       .start_in   (start_in_3_41),
       .op_in      (op_in_3_41),
       .pivot_in   (pivot_in_3_41),
       .start_out  (start_out_3_41),
       .data_out   (data_out_3_41),
       .op_out     (op_out_3_41),
       .pivot_out  (pivot_out_3_41),
       .r          (r_3_41)
     );

  // row 3, col 42

     reg start_in_3_42;
     wire start_out_3_42;

     reg [1:0] op_in_3_42;
     wire [1:0] op_out_3_42;

     wire r_3_42;

     reg data_in_3_42;
     wire data_out_3_42;

     reg pivot_in_3_42;
     wire pivot_out_3_42;

     always @(posedge clk) begin
         op_in_3_42 <= op_out_3_41;
         pivot_in_3_42 <= pivot_out_3_41;
         start_in_3_42 <= start_out_3_41;
     end

     always @(posedge clk) begin
         data_in_3_42 <= data_out_2_42;
     end
  
     processor_AB AB_3_42 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_42),
       .start_in   (start_in_3_42),
       .op_in      (op_in_3_42),
       .pivot_in   (pivot_in_3_42),
       .start_out  (start_out_3_42),
       .data_out   (data_out_3_42),
       .op_out     (op_out_3_42),
       .pivot_out  (pivot_out_3_42),
       .r          (r_3_42)
     );

  // row 3, col 43

     reg start_in_3_43;
     wire start_out_3_43;

     reg [1:0] op_in_3_43;
     wire [1:0] op_out_3_43;

     wire r_3_43;

     reg data_in_3_43;
     wire data_out_3_43;

     reg pivot_in_3_43;
     wire pivot_out_3_43;

     always @(posedge clk) begin
         op_in_3_43 <= op_out_3_42;
         pivot_in_3_43 <= pivot_out_3_42;
         start_in_3_43 <= start_out_3_42;
     end

     always @(posedge clk) begin
         data_in_3_43 <= data_out_2_43;
     end
  
     processor_AB AB_3_43 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_43),
       .start_in   (start_in_3_43),
       .op_in      (op_in_3_43),
       .pivot_in   (pivot_in_3_43),
       .start_out  (start_out_3_43),
       .data_out   (data_out_3_43),
       .op_out     (op_out_3_43),
       .pivot_out  (pivot_out_3_43),
       .r          (r_3_43)
     );

  // row 3, col 44

     reg start_in_3_44;
     wire start_out_3_44;

     reg [1:0] op_in_3_44;
     wire [1:0] op_out_3_44;

     wire r_3_44;

     reg data_in_3_44;
     wire data_out_3_44;

     reg pivot_in_3_44;
     wire pivot_out_3_44;

     always @(posedge clk) begin
         op_in_3_44 <= op_out_3_43;
         pivot_in_3_44 <= pivot_out_3_43;
         start_in_3_44 <= start_out_3_43;
     end

     always @(posedge clk) begin
         data_in_3_44 <= data_out_2_44;
     end
  
     processor_AB AB_3_44 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_44),
       .start_in   (start_in_3_44),
       .op_in      (op_in_3_44),
       .pivot_in   (pivot_in_3_44),
       .start_out  (start_out_3_44),
       .data_out   (data_out_3_44),
       .op_out     (op_out_3_44),
       .pivot_out  (pivot_out_3_44),
       .r          (r_3_44)
     );

  // row 3, col 45

     reg start_in_3_45;
     wire start_out_3_45;

     reg [1:0] op_in_3_45;
     wire [1:0] op_out_3_45;

     wire r_3_45;

     reg data_in_3_45;
     wire data_out_3_45;

     reg pivot_in_3_45;
     wire pivot_out_3_45;

     always @(posedge clk) begin
         op_in_3_45 <= op_out_3_44;
         pivot_in_3_45 <= pivot_out_3_44;
         start_in_3_45 <= start_out_3_44;
     end

     always @(posedge clk) begin
         data_in_3_45 <= data_out_2_45;
     end
  
     processor_AB AB_3_45 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_45),
       .start_in   (start_in_3_45),
       .op_in      (op_in_3_45),
       .pivot_in   (pivot_in_3_45),
       .start_out  (start_out_3_45),
       .data_out   (data_out_3_45),
       .op_out     (op_out_3_45),
       .pivot_out  (pivot_out_3_45),
       .r          (r_3_45)
     );

  // row 3, col 46

     reg start_in_3_46;
     wire start_out_3_46;

     reg [1:0] op_in_3_46;
     wire [1:0] op_out_3_46;

     wire r_3_46;

     reg data_in_3_46;
     wire data_out_3_46;

     reg pivot_in_3_46;
     wire pivot_out_3_46;

     always @(posedge clk) begin
         op_in_3_46 <= op_out_3_45;
         pivot_in_3_46 <= pivot_out_3_45;
         start_in_3_46 <= start_out_3_45;
     end

     always @(posedge clk) begin
         data_in_3_46 <= data_out_2_46;
     end
  
     processor_AB AB_3_46 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_46),
       .start_in   (start_in_3_46),
       .op_in      (op_in_3_46),
       .pivot_in   (pivot_in_3_46),
       .start_out  (start_out_3_46),
       .data_out   (data_out_3_46),
       .op_out     (op_out_3_46),
       .pivot_out  (pivot_out_3_46),
       .r          (r_3_46)
     );

  // row 3, col 47

     reg start_in_3_47;
     wire start_out_3_47;

     reg [1:0] op_in_3_47;
     wire [1:0] op_out_3_47;

     wire r_3_47;

     reg data_in_3_47;
     wire data_out_3_47;

     reg pivot_in_3_47;
     wire pivot_out_3_47;

     always @(posedge clk) begin
         op_in_3_47 <= op_out_3_46;
         pivot_in_3_47 <= pivot_out_3_46;
         start_in_3_47 <= start_out_3_46;
     end

     always @(posedge clk) begin
         data_in_3_47 <= data_out_2_47;
     end
  
     processor_AB AB_3_47 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_47),
       .start_in   (start_in_3_47),
       .op_in      (op_in_3_47),
       .pivot_in   (pivot_in_3_47),
       .start_out  (start_out_3_47),
       .data_out   (data_out_3_47),
       .op_out     (op_out_3_47),
       .pivot_out  (pivot_out_3_47),
       .r          (r_3_47)
     );

  // row 3, col 48

     reg start_in_3_48;
     wire start_out_3_48;

     reg [1:0] op_in_3_48;
     wire [1:0] op_out_3_48;

     wire r_3_48;

     reg data_in_3_48;
     wire data_out_3_48;

     reg pivot_in_3_48;
     wire pivot_out_3_48;

     always @(posedge clk) begin
         op_in_3_48 <= op_out_3_47;
         pivot_in_3_48 <= pivot_out_3_47;
         start_in_3_48 <= start_out_3_47;
     end

     always @(posedge clk) begin
         data_in_3_48 <= data_out_2_48;
     end
  
     processor_AB AB_3_48 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_48),
       .start_in   (start_in_3_48),
       .op_in      (op_in_3_48),
       .pivot_in   (pivot_in_3_48),
       .start_out  (start_out_3_48),
       .data_out   (data_out_3_48),
       .op_out     (op_out_3_48),
       .pivot_out  (pivot_out_3_48),
       .r          (r_3_48)
     );

  // row 3, col 49

     reg start_in_3_49;
     wire start_out_3_49;

     reg [1:0] op_in_3_49;
     wire [1:0] op_out_3_49;

     wire r_3_49;

     reg data_in_3_49;
     wire data_out_3_49;

     reg pivot_in_3_49;
     wire pivot_out_3_49;

     always @(posedge clk) begin
         op_in_3_49 <= op_out_3_48;
         pivot_in_3_49 <= pivot_out_3_48;
         start_in_3_49 <= start_out_3_48;
     end

     always @(posedge clk) begin
         data_in_3_49 <= data_out_2_49;
     end
  
     processor_AB AB_3_49 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_49),
       .start_in   (start_in_3_49),
       .op_in      (op_in_3_49),
       .pivot_in   (pivot_in_3_49),
       .start_out  (start_out_3_49),
       .data_out   (data_out_3_49),
       .op_out     (op_out_3_49),
       .pivot_out  (pivot_out_3_49),
       .r          (r_3_49)
     );

  // row 3, col 50

     reg start_in_3_50;
     wire start_out_3_50;

     reg [1:0] op_in_3_50;
     wire [1:0] op_out_3_50;

     wire r_3_50;

     reg data_in_3_50;
     wire data_out_3_50;

     reg pivot_in_3_50;
     wire pivot_out_3_50;

     always @(posedge clk) begin
         op_in_3_50 <= op_out_3_49;
         pivot_in_3_50 <= pivot_out_3_49;
         start_in_3_50 <= start_out_3_49;
     end

     always @(posedge clk) begin
         data_in_3_50 <= data_out_2_50;
     end
  
     processor_AB AB_3_50 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_50),
       .start_in   (start_in_3_50),
       .op_in      (op_in_3_50),
       .pivot_in   (pivot_in_3_50),
       .start_out  (start_out_3_50),
       .data_out   (data_out_3_50),
       .op_out     (op_out_3_50),
       .pivot_out  (pivot_out_3_50),
       .r          (r_3_50)
     );

  // row 3, col 51

     reg start_in_3_51;
     wire start_out_3_51;

     reg [1:0] op_in_3_51;
     wire [1:0] op_out_3_51;

     wire r_3_51;

     reg data_in_3_51;
     wire data_out_3_51;

     reg pivot_in_3_51;
     wire pivot_out_3_51;

     always @(posedge clk) begin
         op_in_3_51 <= op_out_3_50;
         pivot_in_3_51 <= pivot_out_3_50;
         start_in_3_51 <= start_out_3_50;
     end

     always @(posedge clk) begin
         data_in_3_51 <= data_out_2_51;
     end
  
     processor_AB AB_3_51 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_51),
       .start_in   (start_in_3_51),
       .op_in      (op_in_3_51),
       .pivot_in   (pivot_in_3_51),
       .start_out  (start_out_3_51),
       .data_out   (data_out_3_51),
       .op_out     (op_out_3_51),
       .pivot_out  (pivot_out_3_51),
       .r          (r_3_51)
     );

  // row 3, col 52

     reg start_in_3_52;
     wire start_out_3_52;

     reg [1:0] op_in_3_52;
     wire [1:0] op_out_3_52;

     wire r_3_52;

     reg data_in_3_52;
     wire data_out_3_52;

     reg pivot_in_3_52;
     wire pivot_out_3_52;

     always @(posedge clk) begin
         op_in_3_52 <= op_out_3_51;
         pivot_in_3_52 <= pivot_out_3_51;
         start_in_3_52 <= start_out_3_51;
     end

     always @(posedge clk) begin
         data_in_3_52 <= data_out_2_52;
     end
  
     processor_AB AB_3_52 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_52),
       .start_in   (start_in_3_52),
       .op_in      (op_in_3_52),
       .pivot_in   (pivot_in_3_52),
       .start_out  (start_out_3_52),
       .data_out   (data_out_3_52),
       .op_out     (op_out_3_52),
       .pivot_out  (pivot_out_3_52),
       .r          (r_3_52)
     );

  // row 3, col 53

     reg start_in_3_53;
     wire start_out_3_53;

     reg [1:0] op_in_3_53;
     wire [1:0] op_out_3_53;

     wire r_3_53;

     reg data_in_3_53;
     wire data_out_3_53;

     reg pivot_in_3_53;
     wire pivot_out_3_53;

     always @(posedge clk) begin
         op_in_3_53 <= op_out_3_52;
         pivot_in_3_53 <= pivot_out_3_52;
         start_in_3_53 <= start_out_3_52;
     end

     always @(posedge clk) begin
         data_in_3_53 <= data_out_2_53;
     end
  
     processor_AB AB_3_53 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_53),
       .start_in   (start_in_3_53),
       .op_in      (op_in_3_53),
       .pivot_in   (pivot_in_3_53),
       .start_out  (start_out_3_53),
       .data_out   (data_out_3_53),
       .op_out     (op_out_3_53),
       .pivot_out  (pivot_out_3_53),
       .r          (r_3_53)
     );

  // row 3, col 54

     reg start_in_3_54;
     wire start_out_3_54;

     reg [1:0] op_in_3_54;
     wire [1:0] op_out_3_54;

     wire r_3_54;

     reg data_in_3_54;
     wire data_out_3_54;

     reg pivot_in_3_54;
     wire pivot_out_3_54;

     always @(posedge clk) begin
         op_in_3_54 <= op_out_3_53;
         pivot_in_3_54 <= pivot_out_3_53;
         start_in_3_54 <= start_out_3_53;
     end

     always @(posedge clk) begin
         data_in_3_54 <= data_out_2_54;
     end
  
     processor_AB AB_3_54 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_54),
       .start_in   (start_in_3_54),
       .op_in      (op_in_3_54),
       .pivot_in   (pivot_in_3_54),
       .start_out  (start_out_3_54),
       .data_out   (data_out_3_54),
       .op_out     (op_out_3_54),
       .pivot_out  (pivot_out_3_54),
       .r          (r_3_54)
     );

  // row 3, col 55

     reg start_in_3_55;
     wire start_out_3_55;

     reg [1:0] op_in_3_55;
     wire [1:0] op_out_3_55;

     wire r_3_55;

     reg data_in_3_55;
     wire data_out_3_55;

     reg pivot_in_3_55;
     wire pivot_out_3_55;

     always @(posedge clk) begin
         op_in_3_55 <= op_out_3_54;
         pivot_in_3_55 <= pivot_out_3_54;
         start_in_3_55 <= start_out_3_54;
     end

     always @(posedge clk) begin
         data_in_3_55 <= data_out_2_55;
     end
  
     processor_AB AB_3_55 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_55),
       .start_in   (start_in_3_55),
       .op_in      (op_in_3_55),
       .pivot_in   (pivot_in_3_55),
       .start_out  (start_out_3_55),
       .data_out   (data_out_3_55),
       .op_out     (op_out_3_55),
       .pivot_out  (pivot_out_3_55),
       .r          (r_3_55)
     );

  // row 3, col 56

     reg start_in_3_56;
     wire start_out_3_56;

     reg [1:0] op_in_3_56;
     wire [1:0] op_out_3_56;

     wire r_3_56;

     reg data_in_3_56;
     wire data_out_3_56;

     reg pivot_in_3_56;
     wire pivot_out_3_56;

     always @(posedge clk) begin
         op_in_3_56 <= op_out_3_55;
         pivot_in_3_56 <= pivot_out_3_55;
         start_in_3_56 <= start_out_3_55;
     end

     always @(posedge clk) begin
         data_in_3_56 <= data_out_2_56;
     end
  
     processor_AB AB_3_56 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_56),
       .start_in   (start_in_3_56),
       .op_in      (op_in_3_56),
       .pivot_in   (pivot_in_3_56),
       .start_out  (start_out_3_56),
       .data_out   (data_out_3_56),
       .op_out     (op_out_3_56),
       .pivot_out  (pivot_out_3_56),
       .r          (r_3_56)
     );

  // row 3, col 57

     reg start_in_3_57;
     wire start_out_3_57;

     reg [1:0] op_in_3_57;
     wire [1:0] op_out_3_57;

     wire r_3_57;

     reg data_in_3_57;
     wire data_out_3_57;

     reg pivot_in_3_57;
     wire pivot_out_3_57;

     always @(posedge clk) begin
         op_in_3_57 <= op_out_3_56;
         pivot_in_3_57 <= pivot_out_3_56;
         start_in_3_57 <= start_out_3_56;
     end

     always @(posedge clk) begin
         data_in_3_57 <= data_out_2_57;
     end
  
     processor_AB AB_3_57 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_57),
       .start_in   (start_in_3_57),
       .op_in      (op_in_3_57),
       .pivot_in   (pivot_in_3_57),
       .start_out  (start_out_3_57),
       .data_out   (data_out_3_57),
       .op_out     (op_out_3_57),
       .pivot_out  (pivot_out_3_57),
       .r          (r_3_57)
     );

  // row 3, col 58

     reg start_in_3_58;
     wire start_out_3_58;

     reg [1:0] op_in_3_58;
     wire [1:0] op_out_3_58;

     wire r_3_58;

     reg data_in_3_58;
     wire data_out_3_58;

     reg pivot_in_3_58;
     wire pivot_out_3_58;

     always @(posedge clk) begin
         op_in_3_58 <= op_out_3_57;
         pivot_in_3_58 <= pivot_out_3_57;
         start_in_3_58 <= start_out_3_57;
     end

     always @(posedge clk) begin
         data_in_3_58 <= data_out_2_58;
     end
  
     processor_AB AB_3_58 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_58),
       .start_in   (start_in_3_58),
       .op_in      (op_in_3_58),
       .pivot_in   (pivot_in_3_58),
       .start_out  (start_out_3_58),
       .data_out   (data_out_3_58),
       .op_out     (op_out_3_58),
       .pivot_out  (pivot_out_3_58),
       .r          (r_3_58)
     );

  // row 3, col 59

     reg start_in_3_59;
     wire start_out_3_59;

     reg [1:0] op_in_3_59;
     wire [1:0] op_out_3_59;

     wire r_3_59;

     reg data_in_3_59;
     wire data_out_3_59;

     reg pivot_in_3_59;
     wire pivot_out_3_59;

     always @(posedge clk) begin
         op_in_3_59 <= op_out_3_58;
         pivot_in_3_59 <= pivot_out_3_58;
         start_in_3_59 <= start_out_3_58;
     end

     always @(posedge clk) begin
         data_in_3_59 <= data_out_2_59;
     end
  
     processor_AB AB_3_59 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_59),
       .start_in   (start_in_3_59),
       .op_in      (op_in_3_59),
       .pivot_in   (pivot_in_3_59),
       .start_out  (start_out_3_59),
       .data_out   (data_out_3_59),
       .op_out     (op_out_3_59),
       .pivot_out  (pivot_out_3_59),
       .r          (r_3_59)
     );

  // row 3, col 60

     reg start_in_3_60;
     wire start_out_3_60;

     reg [1:0] op_in_3_60;
     wire [1:0] op_out_3_60;

     wire r_3_60;

     reg data_in_3_60;
     wire data_out_3_60;

     reg pivot_in_3_60;
     wire pivot_out_3_60;

     always @(posedge clk) begin
         op_in_3_60 <= op_out_3_59;
         pivot_in_3_60 <= pivot_out_3_59;
         start_in_3_60 <= start_out_3_59;
     end

     always @(posedge clk) begin
         data_in_3_60 <= data_out_2_60;
     end
  
     processor_AB AB_3_60 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_60),
       .start_in   (start_in_3_60),
       .op_in      (op_in_3_60),
       .pivot_in   (pivot_in_3_60),
       .start_out  (start_out_3_60),
       .data_out   (data_out_3_60),
       .op_out     (op_out_3_60),
       .pivot_out  (pivot_out_3_60),
       .r          (r_3_60)
     );

  // row 3, col 61

     reg start_in_3_61;
     wire start_out_3_61;

     reg [1:0] op_in_3_61;
     wire [1:0] op_out_3_61;

     wire r_3_61;

     reg data_in_3_61;
     wire data_out_3_61;

     reg pivot_in_3_61;
     wire pivot_out_3_61;

     always @(posedge clk) begin
         op_in_3_61 <= op_out_3_60;
         pivot_in_3_61 <= pivot_out_3_60;
         start_in_3_61 <= start_out_3_60;
     end

     always @(posedge clk) begin
         data_in_3_61 <= data_out_2_61;
     end
  
     processor_AB AB_3_61 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_61),
       .start_in   (start_in_3_61),
       .op_in      (op_in_3_61),
       .pivot_in   (pivot_in_3_61),
       .start_out  (start_out_3_61),
       .data_out   (data_out_3_61),
       .op_out     (op_out_3_61),
       .pivot_out  (pivot_out_3_61),
       .r          (r_3_61)
     );

  // row 3, col 62

     reg start_in_3_62;
     wire start_out_3_62;

     reg [1:0] op_in_3_62;
     wire [1:0] op_out_3_62;

     wire r_3_62;

     reg data_in_3_62;
     wire data_out_3_62;

     reg pivot_in_3_62;
     wire pivot_out_3_62;

     always @(posedge clk) begin
         op_in_3_62 <= op_out_3_61;
         pivot_in_3_62 <= pivot_out_3_61;
         start_in_3_62 <= start_out_3_61;
     end

     always @(posedge clk) begin
         data_in_3_62 <= data_out_2_62;
     end
  
     processor_AB AB_3_62 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_62),
       .start_in   (start_in_3_62),
       .op_in      (op_in_3_62),
       .pivot_in   (pivot_in_3_62),
       .start_out  (start_out_3_62),
       .data_out   (data_out_3_62),
       .op_out     (op_out_3_62),
       .pivot_out  (pivot_out_3_62),
       .r          (r_3_62)
     );

  // row 3, col 63

     reg start_in_3_63;
     wire start_out_3_63;

     reg [1:0] op_in_3_63;
     wire [1:0] op_out_3_63;

     wire r_3_63;

     reg data_in_3_63;
     wire data_out_3_63;

     reg pivot_in_3_63;
     wire pivot_out_3_63;

     always @(posedge clk) begin
         op_in_3_63 <= op_out_3_62;
         pivot_in_3_63 <= pivot_out_3_62;
         start_in_3_63 <= start_out_3_62;
     end

     always @(posedge clk) begin
         data_in_3_63 <= data_out_2_63;
     end
  
     processor_AB AB_3_63 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_63),
       .start_in   (start_in_3_63),
       .op_in      (op_in_3_63),
       .pivot_in   (pivot_in_3_63),
       .start_out  (start_out_3_63),
       .data_out   (data_out_3_63),
       .op_out     (op_out_3_63),
       .pivot_out  (pivot_out_3_63),
       .r          (r_3_63)
     );

  // row 3, col 64

     reg start_in_3_64;
     wire start_out_3_64;

     reg [1:0] op_in_3_64;
     wire [1:0] op_out_3_64;

     wire r_3_64;

     reg data_in_3_64;
     wire data_out_3_64;

     reg pivot_in_3_64;
     wire pivot_out_3_64;

     always @(posedge clk) begin
         op_in_3_64 <= op_out_3_63;
         pivot_in_3_64 <= pivot_out_3_63;
         start_in_3_64 <= start_out_3_63;
     end

     always @(posedge clk) begin
         data_in_3_64 <= data_out_2_64;
     end
  
     processor_AB AB_3_64 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_64),
       .start_in   (start_in_3_64),
       .op_in      (op_in_3_64),
       .pivot_in   (pivot_in_3_64),
       .start_out  (start_out_3_64),
       .data_out   (data_out_3_64),
       .op_out     (op_out_3_64),
       .pivot_out  (pivot_out_3_64),
       .r          (r_3_64)
     );

  // row 3, col 65

     reg start_in_3_65;
     wire start_out_3_65;

     reg [1:0] op_in_3_65;
     wire [1:0] op_out_3_65;

     wire r_3_65;

     reg data_in_3_65;
     wire data_out_3_65;

     reg pivot_in_3_65;
     wire pivot_out_3_65;

     always @(posedge clk) begin
         op_in_3_65 <= op_out_3_64;
         pivot_in_3_65 <= pivot_out_3_64;
         start_in_3_65 <= start_out_3_64;
     end

     always @(posedge clk) begin
         data_in_3_65 <= data_out_2_65;
     end
  
     processor_AB AB_3_65 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_65),
       .start_in   (start_in_3_65),
       .op_in      (op_in_3_65),
       .pivot_in   (pivot_in_3_65),
       .start_out  (start_out_3_65),
       .data_out   (data_out_3_65),
       .op_out     (op_out_3_65),
       .pivot_out  (pivot_out_3_65),
       .r          (r_3_65)
     );

  // row 3, col 66

     reg start_in_3_66;
     wire start_out_3_66;

     reg [1:0] op_in_3_66;
     wire [1:0] op_out_3_66;

     wire r_3_66;

     reg data_in_3_66;
     wire data_out_3_66;

     reg pivot_in_3_66;
     wire pivot_out_3_66;

     always @(posedge clk) begin
         op_in_3_66 <= op_out_3_65;
         pivot_in_3_66 <= pivot_out_3_65;
         start_in_3_66 <= start_out_3_65;
     end

     always @(posedge clk) begin
         data_in_3_66 <= data_out_2_66;
     end
  
     processor_AB AB_3_66 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_66),
       .start_in   (start_in_3_66),
       .op_in      (op_in_3_66),
       .pivot_in   (pivot_in_3_66),
       .start_out  (start_out_3_66),
       .data_out   (data_out_3_66),
       .op_out     (op_out_3_66),
       .pivot_out  (pivot_out_3_66),
       .r          (r_3_66)
     );

  // row 3, col 67

     reg start_in_3_67;
     wire start_out_3_67;

     reg [1:0] op_in_3_67;
     wire [1:0] op_out_3_67;

     wire r_3_67;

     reg data_in_3_67;
     wire data_out_3_67;

     reg pivot_in_3_67;
     wire pivot_out_3_67;

     always @(posedge clk) begin
         op_in_3_67 <= op_out_3_66;
         pivot_in_3_67 <= pivot_out_3_66;
         start_in_3_67 <= start_out_3_66;
     end

     always @(posedge clk) begin
         data_in_3_67 <= data_out_2_67;
     end
  
     processor_AB AB_3_67 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_67),
       .start_in   (start_in_3_67),
       .op_in      (op_in_3_67),
       .pivot_in   (pivot_in_3_67),
       .start_out  (start_out_3_67),
       .data_out   (data_out_3_67),
       .op_out     (op_out_3_67),
       .pivot_out  (pivot_out_3_67),
       .r          (r_3_67)
     );

  // row 3, col 68

     reg start_in_3_68;
     wire start_out_3_68;

     reg [1:0] op_in_3_68;
     wire [1:0] op_out_3_68;

     wire r_3_68;

     reg data_in_3_68;
     wire data_out_3_68;

     reg pivot_in_3_68;
     wire pivot_out_3_68;

     always @(posedge clk) begin
         op_in_3_68 <= op_out_3_67;
         pivot_in_3_68 <= pivot_out_3_67;
         start_in_3_68 <= start_out_3_67;
     end

     always @(posedge clk) begin
         data_in_3_68 <= data_out_2_68;
     end
  
     processor_AB AB_3_68 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_68),
       .start_in   (start_in_3_68),
       .op_in      (op_in_3_68),
       .pivot_in   (pivot_in_3_68),
       .start_out  (start_out_3_68),
       .data_out   (data_out_3_68),
       .op_out     (op_out_3_68),
       .pivot_out  (pivot_out_3_68),
       .r          (r_3_68)
     );

  // row 3, col 69

     reg start_in_3_69;
     wire start_out_3_69;

     reg [1:0] op_in_3_69;
     wire [1:0] op_out_3_69;

     wire r_3_69;

     reg data_in_3_69;
     wire data_out_3_69;

     reg pivot_in_3_69;
     wire pivot_out_3_69;

     always @(posedge clk) begin
         op_in_3_69 <= op_out_3_68;
         pivot_in_3_69 <= pivot_out_3_68;
         start_in_3_69 <= start_out_3_68;
     end

     always @(posedge clk) begin
         data_in_3_69 <= data_out_2_69;
     end
  
     processor_AB AB_3_69 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_69),
       .start_in   (start_in_3_69),
       .op_in      (op_in_3_69),
       .pivot_in   (pivot_in_3_69),
       .start_out  (start_out_3_69),
       .data_out   (data_out_3_69),
       .op_out     (op_out_3_69),
       .pivot_out  (pivot_out_3_69),
       .r          (r_3_69)
     );

  // row 3, col 70

     reg start_in_3_70;
     wire start_out_3_70;

     reg [1:0] op_in_3_70;
     wire [1:0] op_out_3_70;

     wire r_3_70;

     reg data_in_3_70;
     wire data_out_3_70;

     reg pivot_in_3_70;
     wire pivot_out_3_70;

     always @(posedge clk) begin
         op_in_3_70 <= op_out_3_69;
         pivot_in_3_70 <= pivot_out_3_69;
         start_in_3_70 <= start_out_3_69;
     end

     always @(posedge clk) begin
         data_in_3_70 <= data_out_2_70;
     end
  
     processor_AB AB_3_70 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_70),
       .start_in   (start_in_3_70),
       .op_in      (op_in_3_70),
       .pivot_in   (pivot_in_3_70),
       .start_out  (start_out_3_70),
       .data_out   (data_out_3_70),
       .op_out     (op_out_3_70),
       .pivot_out  (pivot_out_3_70),
       .r          (r_3_70)
     );

  // row 3, col 71

     reg start_in_3_71;
     wire start_out_3_71;

     reg [1:0] op_in_3_71;
     wire [1:0] op_out_3_71;

     wire r_3_71;

     reg data_in_3_71;
     wire data_out_3_71;

     reg pivot_in_3_71;
     wire pivot_out_3_71;

     always @(posedge clk) begin
         op_in_3_71 <= op_out_3_70;
         pivot_in_3_71 <= pivot_out_3_70;
         start_in_3_71 <= start_out_3_70;
     end

     always @(posedge clk) begin
         data_in_3_71 <= data_out_2_71;
     end
  
     processor_AB AB_3_71 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_71),
       .start_in   (start_in_3_71),
       .op_in      (op_in_3_71),
       .pivot_in   (pivot_in_3_71),
       .start_out  (start_out_3_71),
       .data_out   (data_out_3_71),
       .op_out     (op_out_3_71),
       .pivot_out  (pivot_out_3_71),
       .r          (r_3_71)
     );

  // row 3, col 72

     reg start_in_3_72;
     wire start_out_3_72;

     reg [1:0] op_in_3_72;
     wire [1:0] op_out_3_72;

     wire r_3_72;

     reg data_in_3_72;
     wire data_out_3_72;

     reg pivot_in_3_72;
     wire pivot_out_3_72;

     always @(posedge clk) begin
         op_in_3_72 <= op_out_3_71;
         pivot_in_3_72 <= pivot_out_3_71;
         start_in_3_72 <= start_out_3_71;
     end

     always @(posedge clk) begin
         data_in_3_72 <= data_out_2_72;
     end
  
     processor_AB AB_3_72 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_72),
       .start_in   (start_in_3_72),
       .op_in      (op_in_3_72),
       .pivot_in   (pivot_in_3_72),
       .start_out  (start_out_3_72),
       .data_out   (data_out_3_72),
       .op_out     (op_out_3_72),
       .pivot_out  (pivot_out_3_72),
       .r          (r_3_72)
     );

  // row 3, col 73

     reg start_in_3_73;
     wire start_out_3_73;

     reg [1:0] op_in_3_73;
     wire [1:0] op_out_3_73;

     wire r_3_73;

     reg data_in_3_73;
     wire data_out_3_73;

     reg pivot_in_3_73;
     wire pivot_out_3_73;

     always @(posedge clk) begin
         op_in_3_73 <= op_out_3_72;
         pivot_in_3_73 <= pivot_out_3_72;
         start_in_3_73 <= start_out_3_72;
     end

     always @(posedge clk) begin
         data_in_3_73 <= data_out_2_73;
     end
  
     processor_AB AB_3_73 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_73),
       .start_in   (start_in_3_73),
       .op_in      (op_in_3_73),
       .pivot_in   (pivot_in_3_73),
       .start_out  (start_out_3_73),
       .data_out   (data_out_3_73),
       .op_out     (op_out_3_73),
       .pivot_out  (pivot_out_3_73),
       .r          (r_3_73)
     );

  // row 3, col 74

     reg start_in_3_74;
     wire start_out_3_74;

     reg [1:0] op_in_3_74;
     wire [1:0] op_out_3_74;

     wire r_3_74;

     reg data_in_3_74;
     wire data_out_3_74;

     reg pivot_in_3_74;
     wire pivot_out_3_74;

     always @(posedge clk) begin
         op_in_3_74 <= op_out_3_73;
         pivot_in_3_74 <= pivot_out_3_73;
         start_in_3_74 <= start_out_3_73;
     end

     always @(posedge clk) begin
         data_in_3_74 <= data_out_2_74;
     end
  
     processor_AB AB_3_74 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_74),
       .start_in   (start_in_3_74),
       .op_in      (op_in_3_74),
       .pivot_in   (pivot_in_3_74),
       .start_out  (start_out_3_74),
       .data_out   (data_out_3_74),
       .op_out     (op_out_3_74),
       .pivot_out  (pivot_out_3_74),
       .r          (r_3_74)
     );

  // row 3, col 75

     reg start_in_3_75;
     wire start_out_3_75;

     reg [1:0] op_in_3_75;
     wire [1:0] op_out_3_75;

     wire r_3_75;

     reg data_in_3_75;
     wire data_out_3_75;

     reg pivot_in_3_75;
     wire pivot_out_3_75;

     always @(posedge clk) begin
         op_in_3_75 <= op_out_3_74;
         pivot_in_3_75 <= pivot_out_3_74;
         start_in_3_75 <= start_out_3_74;
     end

     always @(posedge clk) begin
         data_in_3_75 <= data_out_2_75;
     end
  
     processor_AB AB_3_75 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_75),
       .start_in   (start_in_3_75),
       .op_in      (op_in_3_75),
       .pivot_in   (pivot_in_3_75),
       .start_out  (start_out_3_75),
       .data_out   (data_out_3_75),
       .op_out     (op_out_3_75),
       .pivot_out  (pivot_out_3_75),
       .r          (r_3_75)
     );

  // row 3, col 76

     reg start_in_3_76;
     wire start_out_3_76;

     reg [1:0] op_in_3_76;
     wire [1:0] op_out_3_76;

     wire r_3_76;

     reg data_in_3_76;
     wire data_out_3_76;

     reg pivot_in_3_76;
     wire pivot_out_3_76;

     always @(posedge clk) begin
         op_in_3_76 <= op_out_3_75;
         pivot_in_3_76 <= pivot_out_3_75;
         start_in_3_76 <= start_out_3_75;
     end

     always @(posedge clk) begin
         data_in_3_76 <= data_out_2_76;
     end
  
     processor_AB AB_3_76 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_76),
       .start_in   (start_in_3_76),
       .op_in      (op_in_3_76),
       .pivot_in   (pivot_in_3_76),
       .start_out  (start_out_3_76),
       .data_out   (data_out_3_76),
       .op_out     (op_out_3_76),
       .pivot_out  (pivot_out_3_76),
       .r          (r_3_76)
     );

  // row 3, col 77

     reg start_in_3_77;
     wire start_out_3_77;

     reg [1:0] op_in_3_77;
     wire [1:0] op_out_3_77;

     wire r_3_77;

     reg data_in_3_77;
     wire data_out_3_77;

     reg pivot_in_3_77;
     wire pivot_out_3_77;

     always @(posedge clk) begin
         op_in_3_77 <= op_out_3_76;
         pivot_in_3_77 <= pivot_out_3_76;
         start_in_3_77 <= start_out_3_76;
     end

     always @(posedge clk) begin
         data_in_3_77 <= data_out_2_77;
     end
  
     processor_AB AB_3_77 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_77),
       .start_in   (start_in_3_77),
       .op_in      (op_in_3_77),
       .pivot_in   (pivot_in_3_77),
       .start_out  (start_out_3_77),
       .data_out   (data_out_3_77),
       .op_out     (op_out_3_77),
       .pivot_out  (pivot_out_3_77),
       .r          (r_3_77)
     );

  // row 3, col 78

     reg start_in_3_78;
     wire start_out_3_78;

     reg [1:0] op_in_3_78;
     wire [1:0] op_out_3_78;

     wire r_3_78;

     reg data_in_3_78;
     wire data_out_3_78;

     reg pivot_in_3_78;
     wire pivot_out_3_78;

     always @(posedge clk) begin
         op_in_3_78 <= op_out_3_77;
         pivot_in_3_78 <= pivot_out_3_77;
         start_in_3_78 <= start_out_3_77;
     end

     always @(posedge clk) begin
         data_in_3_78 <= data_out_2_78;
     end
  
     processor_AB AB_3_78 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_78),
       .start_in   (start_in_3_78),
       .op_in      (op_in_3_78),
       .pivot_in   (pivot_in_3_78),
       .start_out  (start_out_3_78),
       .data_out   (data_out_3_78),
       .op_out     (op_out_3_78),
       .pivot_out  (pivot_out_3_78),
       .r          (r_3_78)
     );

  // row 3, col 79

     reg start_in_3_79;
     wire start_out_3_79;

     reg [1:0] op_in_3_79;
     wire [1:0] op_out_3_79;

     wire r_3_79;

     reg data_in_3_79;
     wire data_out_3_79;

     reg pivot_in_3_79;
     wire pivot_out_3_79;

     always @(posedge clk) begin
         op_in_3_79 <= op_out_3_78;
         pivot_in_3_79 <= pivot_out_3_78;
         start_in_3_79 <= start_out_3_78;
     end

     always @(posedge clk) begin
         data_in_3_79 <= data_out_2_79;
     end
  
     processor_AB AB_3_79 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_79),
       .start_in   (start_in_3_79),
       .op_in      (op_in_3_79),
       .pivot_in   (pivot_in_3_79),
       .start_out  (start_out_3_79),
       .data_out   (data_out_3_79),
       .op_out     (op_out_3_79),
       .pivot_out  (pivot_out_3_79),
       .r          (r_3_79)
     );

  // row 3, col 80

     reg start_in_3_80;
     wire start_out_3_80;

     reg [1:0] op_in_3_80;
     wire [1:0] op_out_3_80;

     wire r_3_80;

     reg data_in_3_80;
     wire data_out_3_80;

     reg pivot_in_3_80;
     wire pivot_out_3_80;

     always @(posedge clk) begin
         op_in_3_80 <= op_out_3_79;
         pivot_in_3_80 <= pivot_out_3_79;
         start_in_3_80 <= start_out_3_79;
     end

     always @(posedge clk) begin
         data_in_3_80 <= data_out_2_80;
     end
  
     processor_AB AB_3_80 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_80),
       .start_in   (start_in_3_80),
       .op_in      (op_in_3_80),
       .pivot_in   (pivot_in_3_80),
       .start_out  (start_out_3_80),
       .data_out   (data_out_3_80),
       .op_out     (op_out_3_80),
       .pivot_out  (pivot_out_3_80),
       .r          (r_3_80)
     );

  // row 3, col 81

     reg start_in_3_81;
     wire start_out_3_81;

     reg [1:0] op_in_3_81;
     wire [1:0] op_out_3_81;

     wire r_3_81;

     reg data_in_3_81;
     wire data_out_3_81;

     reg pivot_in_3_81;
     wire pivot_out_3_81;

     always @(posedge clk) begin
         op_in_3_81 <= op_out_3_80;
         pivot_in_3_81 <= pivot_out_3_80;
         start_in_3_81 <= start_out_3_80;
     end

     always @(posedge clk) begin
         data_in_3_81 <= data_out_2_81;
     end
  
     processor_AB AB_3_81 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_81),
       .start_in   (start_in_3_81),
       .op_in      (op_in_3_81),
       .pivot_in   (pivot_in_3_81),
       .start_out  (start_out_3_81),
       .data_out   (data_out_3_81),
       .op_out     (op_out_3_81),
       .pivot_out  (pivot_out_3_81),
       .r          (r_3_81)
     );

  // row 3, col 82

     reg start_in_3_82;
     wire start_out_3_82;

     reg [1:0] op_in_3_82;
     wire [1:0] op_out_3_82;

     wire r_3_82;

     reg data_in_3_82;
     wire data_out_3_82;

     reg pivot_in_3_82;
     wire pivot_out_3_82;

     always @(posedge clk) begin
         op_in_3_82 <= op_out_3_81;
         pivot_in_3_82 <= pivot_out_3_81;
         start_in_3_82 <= start_out_3_81;
     end

     always @(posedge clk) begin
         data_in_3_82 <= data_out_2_82;
     end
  
     processor_AB AB_3_82 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_82),
       .start_in   (start_in_3_82),
       .op_in      (op_in_3_82),
       .pivot_in   (pivot_in_3_82),
       .start_out  (start_out_3_82),
       .data_out   (data_out_3_82),
       .op_out     (op_out_3_82),
       .pivot_out  (pivot_out_3_82),
       .r          (r_3_82)
     );

  // row 3, col 83

     reg start_in_3_83;
     wire start_out_3_83;

     reg [1:0] op_in_3_83;
     wire [1:0] op_out_3_83;

     wire r_3_83;

     reg data_in_3_83;
     wire data_out_3_83;

     reg pivot_in_3_83;
     wire pivot_out_3_83;

     always @(posedge clk) begin
         op_in_3_83 <= op_out_3_82;
         pivot_in_3_83 <= pivot_out_3_82;
         start_in_3_83 <= start_out_3_82;
     end

     always @(posedge clk) begin
         data_in_3_83 <= data_out_2_83;
     end
  
     processor_AB AB_3_83 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_83),
       .start_in   (start_in_3_83),
       .op_in      (op_in_3_83),
       .pivot_in   (pivot_in_3_83),
       .start_out  (start_out_3_83),
       .data_out   (data_out_3_83),
       .op_out     (op_out_3_83),
       .pivot_out  (pivot_out_3_83),
       .r          (r_3_83)
     );

  // row 3, col 84

     reg start_in_3_84;
     wire start_out_3_84;

     reg [1:0] op_in_3_84;
     wire [1:0] op_out_3_84;

     wire r_3_84;

     reg data_in_3_84;
     wire data_out_3_84;

     reg pivot_in_3_84;
     wire pivot_out_3_84;

     always @(posedge clk) begin
         op_in_3_84 <= op_out_3_83;
         pivot_in_3_84 <= pivot_out_3_83;
         start_in_3_84 <= start_out_3_83;
     end

     always @(posedge clk) begin
         data_in_3_84 <= data_out_2_84;
     end
  
     processor_AB AB_3_84 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_84),
       .start_in   (start_in_3_84),
       .op_in      (op_in_3_84),
       .pivot_in   (pivot_in_3_84),
       .start_out  (start_out_3_84),
       .data_out   (data_out_3_84),
       .op_out     (op_out_3_84),
       .pivot_out  (pivot_out_3_84),
       .r          (r_3_84)
     );

  // row 3, col 85

     reg start_in_3_85;
     wire start_out_3_85;

     reg [1:0] op_in_3_85;
     wire [1:0] op_out_3_85;

     wire r_3_85;

     reg data_in_3_85;
     wire data_out_3_85;

     reg pivot_in_3_85;
     wire pivot_out_3_85;

     always @(posedge clk) begin
         op_in_3_85 <= op_out_3_84;
         pivot_in_3_85 <= pivot_out_3_84;
         start_in_3_85 <= start_out_3_84;
     end

     always @(posedge clk) begin
         data_in_3_85 <= data_out_2_85;
     end
  
     processor_AB AB_3_85 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_85),
       .start_in   (start_in_3_85),
       .op_in      (op_in_3_85),
       .pivot_in   (pivot_in_3_85),
       .start_out  (start_out_3_85),
       .data_out   (data_out_3_85),
       .op_out     (op_out_3_85),
       .pivot_out  (pivot_out_3_85),
       .r          (r_3_85)
     );

  // row 3, col 86

     reg start_in_3_86;
     wire start_out_3_86;

     reg [1:0] op_in_3_86;
     wire [1:0] op_out_3_86;

     wire r_3_86;

     reg data_in_3_86;
     wire data_out_3_86;

     reg pivot_in_3_86;
     wire pivot_out_3_86;

     always @(posedge clk) begin
         op_in_3_86 <= op_out_3_85;
         pivot_in_3_86 <= pivot_out_3_85;
         start_in_3_86 <= start_out_3_85;
     end

     always @(posedge clk) begin
         data_in_3_86 <= data_out_2_86;
     end
  
     processor_AB AB_3_86 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_86),
       .start_in   (start_in_3_86),
       .op_in      (op_in_3_86),
       .pivot_in   (pivot_in_3_86),
       .start_out  (start_out_3_86),
       .data_out   (data_out_3_86),
       .op_out     (op_out_3_86),
       .pivot_out  (pivot_out_3_86),
       .r          (r_3_86)
     );

  // row 3, col 87

     reg start_in_3_87;
     wire start_out_3_87;

     reg [1:0] op_in_3_87;
     wire [1:0] op_out_3_87;

     wire r_3_87;

     reg data_in_3_87;
     wire data_out_3_87;

     reg pivot_in_3_87;
     wire pivot_out_3_87;

     always @(posedge clk) begin
         op_in_3_87 <= op_out_3_86;
         pivot_in_3_87 <= pivot_out_3_86;
         start_in_3_87 <= start_out_3_86;
     end

     always @(posedge clk) begin
         data_in_3_87 <= data_out_2_87;
     end
  
     processor_AB AB_3_87 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_87),
       .start_in   (start_in_3_87),
       .op_in      (op_in_3_87),
       .pivot_in   (pivot_in_3_87),
       .start_out  (start_out_3_87),
       .data_out   (data_out_3_87),
       .op_out     (op_out_3_87),
       .pivot_out  (pivot_out_3_87),
       .r          (r_3_87)
     );

  // row 3, col 88

     reg start_in_3_88;
     wire start_out_3_88;

     reg [1:0] op_in_3_88;
     wire [1:0] op_out_3_88;

     wire r_3_88;

     reg data_in_3_88;
     wire data_out_3_88;

     reg pivot_in_3_88;
     wire pivot_out_3_88;

     always @(posedge clk) begin
         op_in_3_88 <= op_out_3_87;
         pivot_in_3_88 <= pivot_out_3_87;
         start_in_3_88 <= start_out_3_87;
     end

     always @(posedge clk) begin
         data_in_3_88 <= data_out_2_88;
     end
  
     processor_AB AB_3_88 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_88),
       .start_in   (start_in_3_88),
       .op_in      (op_in_3_88),
       .pivot_in   (pivot_in_3_88),
       .start_out  (start_out_3_88),
       .data_out   (data_out_3_88),
       .op_out     (op_out_3_88),
       .pivot_out  (pivot_out_3_88),
       .r          (r_3_88)
     );

  // row 3, col 89

     reg start_in_3_89;
     wire start_out_3_89;

     reg [1:0] op_in_3_89;
     wire [1:0] op_out_3_89;

     wire r_3_89;

     reg data_in_3_89;
     wire data_out_3_89;

     reg pivot_in_3_89;
     wire pivot_out_3_89;

     always @(posedge clk) begin
         op_in_3_89 <= op_out_3_88;
         pivot_in_3_89 <= pivot_out_3_88;
         start_in_3_89 <= start_out_3_88;
     end

     always @(posedge clk) begin
         data_in_3_89 <= data_out_2_89;
     end
  
     processor_AB AB_3_89 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_89),
       .start_in   (start_in_3_89),
       .op_in      (op_in_3_89),
       .pivot_in   (pivot_in_3_89),
       .start_out  (start_out_3_89),
       .data_out   (data_out_3_89),
       .op_out     (op_out_3_89),
       .pivot_out  (pivot_out_3_89),
       .r          (r_3_89)
     );

  // row 3, col 90

     reg start_in_3_90;
     wire start_out_3_90;

     reg [1:0] op_in_3_90;
     wire [1:0] op_out_3_90;

     wire r_3_90;

     reg data_in_3_90;
     wire data_out_3_90;

     reg pivot_in_3_90;
     wire pivot_out_3_90;

     always @(posedge clk) begin
         op_in_3_90 <= op_out_3_89;
         pivot_in_3_90 <= pivot_out_3_89;
         start_in_3_90 <= start_out_3_89;
     end

     always @(posedge clk) begin
         data_in_3_90 <= data_out_2_90;
     end
  
     processor_AB AB_3_90 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_90),
       .start_in   (start_in_3_90),
       .op_in      (op_in_3_90),
       .pivot_in   (pivot_in_3_90),
       .start_out  (start_out_3_90),
       .data_out   (data_out_3_90),
       .op_out     (op_out_3_90),
       .pivot_out  (pivot_out_3_90),
       .r          (r_3_90)
     );

  // row 3, col 91

     reg start_in_3_91;
     wire start_out_3_91;

     reg [1:0] op_in_3_91;
     wire [1:0] op_out_3_91;

     wire r_3_91;

     reg data_in_3_91;
     wire data_out_3_91;

     reg pivot_in_3_91;
     wire pivot_out_3_91;

     always @(posedge clk) begin
         op_in_3_91 <= op_out_3_90;
         pivot_in_3_91 <= pivot_out_3_90;
         start_in_3_91 <= start_out_3_90;
     end

     always @(posedge clk) begin
         data_in_3_91 <= data_out_2_91;
     end
  
     processor_AB AB_3_91 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_91),
       .start_in   (start_in_3_91),
       .op_in      (op_in_3_91),
       .pivot_in   (pivot_in_3_91),
       .start_out  (start_out_3_91),
       .data_out   (data_out_3_91),
       .op_out     (op_out_3_91),
       .pivot_out  (pivot_out_3_91),
       .r          (r_3_91)
     );

  // row 3, col 92

     reg start_in_3_92;
     wire start_out_3_92;

     reg [1:0] op_in_3_92;
     wire [1:0] op_out_3_92;

     wire r_3_92;

     reg data_in_3_92;
     wire data_out_3_92;

     reg pivot_in_3_92;
     wire pivot_out_3_92;

     always @(posedge clk) begin
         op_in_3_92 <= op_out_3_91;
         pivot_in_3_92 <= pivot_out_3_91;
         start_in_3_92 <= start_out_3_91;
     end

     always @(posedge clk) begin
         data_in_3_92 <= data_out_2_92;
     end
  
     processor_AB AB_3_92 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_92),
       .start_in   (start_in_3_92),
       .op_in      (op_in_3_92),
       .pivot_in   (pivot_in_3_92),
       .start_out  (start_out_3_92),
       .data_out   (data_out_3_92),
       .op_out     (op_out_3_92),
       .pivot_out  (pivot_out_3_92),
       .r          (r_3_92)
     );

  // row 3, col 93

     reg start_in_3_93;
     wire start_out_3_93;

     reg [1:0] op_in_3_93;
     wire [1:0] op_out_3_93;

     wire r_3_93;

     reg data_in_3_93;
     wire data_out_3_93;

     reg pivot_in_3_93;
     wire pivot_out_3_93;

     always @(posedge clk) begin
         op_in_3_93 <= op_out_3_92;
         pivot_in_3_93 <= pivot_out_3_92;
         start_in_3_93 <= start_out_3_92;
     end

     always @(posedge clk) begin
         data_in_3_93 <= data_out_2_93;
     end
  
     processor_AB AB_3_93 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_93),
       .start_in   (start_in_3_93),
       .op_in      (op_in_3_93),
       .pivot_in   (pivot_in_3_93),
       .start_out  (start_out_3_93),
       .data_out   (data_out_3_93),
       .op_out     (op_out_3_93),
       .pivot_out  (pivot_out_3_93),
       .r          (r_3_93)
     );

  // row 3, col 94

     reg start_in_3_94;
     wire start_out_3_94;

     reg [1:0] op_in_3_94;
     wire [1:0] op_out_3_94;

     wire r_3_94;

     reg data_in_3_94;
     wire data_out_3_94;

     reg pivot_in_3_94;
     wire pivot_out_3_94;

     always @(posedge clk) begin
         op_in_3_94 <= op_out_3_93;
         pivot_in_3_94 <= pivot_out_3_93;
         start_in_3_94 <= start_out_3_93;
     end

     always @(posedge clk) begin
         data_in_3_94 <= data_out_2_94;
     end
  
     processor_AB AB_3_94 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_94),
       .start_in   (start_in_3_94),
       .op_in      (op_in_3_94),
       .pivot_in   (pivot_in_3_94),
       .start_out  (start_out_3_94),
       .data_out   (data_out_3_94),
       .op_out     (op_out_3_94),
       .pivot_out  (pivot_out_3_94),
       .r          (r_3_94)
     );

  // row 3, col 95

     reg start_in_3_95;
     wire start_out_3_95;

     reg [1:0] op_in_3_95;
     wire [1:0] op_out_3_95;

     wire r_3_95;

     reg data_in_3_95;
     wire data_out_3_95;

     reg pivot_in_3_95;
     wire pivot_out_3_95;

     always @(posedge clk) begin
         op_in_3_95 <= op_out_3_94;
         pivot_in_3_95 <= pivot_out_3_94;
         start_in_3_95 <= start_out_3_94;
     end

     always @(posedge clk) begin
         data_in_3_95 <= data_out_2_95;
     end
  
     processor_AB AB_3_95 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_95),
       .start_in   (start_in_3_95),
       .op_in      (op_in_3_95),
       .pivot_in   (pivot_in_3_95),
       .start_out  (start_out_3_95),
       .data_out   (data_out_3_95),
       .op_out     (op_out_3_95),
       .pivot_out  (pivot_out_3_95),
       .r          (r_3_95)
     );

  // row 3, col 96

     reg start_in_3_96;
     wire start_out_3_96;

     reg [1:0] op_in_3_96;
     wire [1:0] op_out_3_96;

     wire r_3_96;

     reg data_in_3_96;
     wire data_out_3_96;

     reg pivot_in_3_96;
     wire pivot_out_3_96;

     always @(posedge clk) begin
         op_in_3_96 <= op_out_3_95;
         pivot_in_3_96 <= pivot_out_3_95;
         start_in_3_96 <= start_out_3_95;
     end

     always @(posedge clk) begin
         data_in_3_96 <= data_out_2_96;
     end
  
     processor_AB AB_3_96 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_96),
       .start_in   (start_in_3_96),
       .op_in      (op_in_3_96),
       .pivot_in   (pivot_in_3_96),
       .start_out  (start_out_3_96),
       .data_out   (data_out_3_96),
       .op_out     (op_out_3_96),
       .pivot_out  (pivot_out_3_96),
       .r          (r_3_96)
     );

  // row 3, col 97

     reg start_in_3_97;
     wire start_out_3_97;

     reg [1:0] op_in_3_97;
     wire [1:0] op_out_3_97;

     wire r_3_97;

     reg data_in_3_97;
     wire data_out_3_97;

     reg pivot_in_3_97;
     wire pivot_out_3_97;

     always @(posedge clk) begin
         op_in_3_97 <= op_out_3_96;
         pivot_in_3_97 <= pivot_out_3_96;
         start_in_3_97 <= start_out_3_96;
     end

     always @(posedge clk) begin
         data_in_3_97 <= data_out_2_97;
     end
  
     processor_AB AB_3_97 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_97),
       .start_in   (start_in_3_97),
       .op_in      (op_in_3_97),
       .pivot_in   (pivot_in_3_97),
       .start_out  (start_out_3_97),
       .data_out   (data_out_3_97),
       .op_out     (op_out_3_97),
       .pivot_out  (pivot_out_3_97),
       .r          (r_3_97)
     );

  // row 3, col 98

     reg start_in_3_98;
     wire start_out_3_98;

     reg [1:0] op_in_3_98;
     wire [1:0] op_out_3_98;

     wire r_3_98;

     reg data_in_3_98;
     wire data_out_3_98;

     reg pivot_in_3_98;
     wire pivot_out_3_98;

     always @(posedge clk) begin
         op_in_3_98 <= op_out_3_97;
         pivot_in_3_98 <= pivot_out_3_97;
         start_in_3_98 <= start_out_3_97;
     end

     always @(posedge clk) begin
         data_in_3_98 <= data_out_2_98;
     end
  
     processor_AB AB_3_98 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_98),
       .start_in   (start_in_3_98),
       .op_in      (op_in_3_98),
       .pivot_in   (pivot_in_3_98),
       .start_out  (start_out_3_98),
       .data_out   (data_out_3_98),
       .op_out     (op_out_3_98),
       .pivot_out  (pivot_out_3_98),
       .r          (r_3_98)
     );

  // row 3, col 99

     reg start_in_3_99;
     wire start_out_3_99;

     reg [1:0] op_in_3_99;
     wire [1:0] op_out_3_99;

     wire r_3_99;

     reg data_in_3_99;
     wire data_out_3_99;

     reg pivot_in_3_99;
     wire pivot_out_3_99;

     always @(posedge clk) begin
         op_in_3_99 <= op_out_3_98;
         pivot_in_3_99 <= pivot_out_3_98;
         start_in_3_99 <= start_out_3_98;
     end

     always @(posedge clk) begin
         data_in_3_99 <= data_out_2_99;
     end
  
     processor_AB AB_3_99 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_99),
       .start_in   (start_in_3_99),
       .op_in      (op_in_3_99),
       .pivot_in   (pivot_in_3_99),
       .start_out  (start_out_3_99),
       .data_out   (data_out_3_99),
       .op_out     (op_out_3_99),
       .pivot_out  (pivot_out_3_99),
       .r          (r_3_99)
     );

  // row 3, col 100

     reg start_in_3_100;
     wire start_out_3_100;

     reg [1:0] op_in_3_100;
     wire [1:0] op_out_3_100;

     wire r_3_100;

     reg data_in_3_100;
     wire data_out_3_100;

     reg pivot_in_3_100;
     wire pivot_out_3_100;

     always @(posedge clk) begin
         op_in_3_100 <= op_out_3_99;
         pivot_in_3_100 <= pivot_out_3_99;
         start_in_3_100 <= start_out_3_99;
     end

     always @(posedge clk) begin
         data_in_3_100 <= data_out_2_100;
     end
  
     processor_AB AB_3_100 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_100),
       .start_in   (start_in_3_100),
       .op_in      (op_in_3_100),
       .pivot_in   (pivot_in_3_100),
       .start_out  (start_out_3_100),
       .data_out   (data_out_3_100),
       .op_out     (op_out_3_100),
       .pivot_out  (pivot_out_3_100),
       .r          (r_3_100)
     );

  /////////////////////////////////////
  // row 4
  // row 4, col 0

     wire start_in_4_0;
     wire start_out_4_0;

     wire [1:0] op_in_4_0;
     wire [1:0] op_out_4_0;

     wire r_4_0;

     reg data_in_4_0;
     wire data_out_4_0;

     wire pivot_in_4_0;
     wire pivout_out_4_0;

     assign op_in_4_0 = mode & start ? 2'b01 : 2'b00;
     assign pivot_in_4_0 = 0;

     assign start_in_4_0 = start_row[4]; 

     always @(posedge clk) begin
         data_in_4_0 <= data_out_3_0;
     end

     processor_AB AB_4_0 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_0),
       .start_in   (start_in_4_0),
       .op_in      (op_in_4_0),
       .pivot_in   (pivot_in_4_0),
       .start_out  (start_out_4_0),
       .data_out   (data_out_4_0),
       .op_out     (op_out_4_0),
       .pivot_out  (pivot_out_4_0),
       .r          (r_4_0)
     );

  // row 4, col 1

     reg start_in_4_1;
     wire start_out_4_1;

     reg [1:0] op_in_4_1;
     wire [1:0] op_out_4_1;

     wire r_4_1;

     reg data_in_4_1;
     wire data_out_4_1;

     reg pivot_in_4_1;
     wire pivot_out_4_1;

     always @(posedge clk) begin
         op_in_4_1 <= op_out_4_0;
         pivot_in_4_1 <= pivot_out_4_0;
         start_in_4_1 <= start_out_4_0;
     end

     always @(posedge clk) begin
         data_in_4_1 <= data_out_3_1;
     end
  
     processor_AB AB_4_1 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_1),
       .start_in   (start_in_4_1),
       .op_in      (op_in_4_1),
       .pivot_in   (pivot_in_4_1),
       .start_out  (start_out_4_1),
       .data_out   (data_out_4_1),
       .op_out     (op_out_4_1),
       .pivot_out  (pivot_out_4_1),
       .r          (r_4_1)
     );

  // row 4, col 2

     reg start_in_4_2;
     wire start_out_4_2;

     reg [1:0] op_in_4_2;
     wire [1:0] op_out_4_2;

     wire r_4_2;

     reg data_in_4_2;
     wire data_out_4_2;

     reg pivot_in_4_2;
     wire pivot_out_4_2;

     always @(posedge clk) begin
         op_in_4_2 <= op_out_4_1;
         pivot_in_4_2 <= pivot_out_4_1;
         start_in_4_2 <= start_out_4_1;
     end

     always @(posedge clk) begin
         data_in_4_2 <= data_out_3_2;
     end
  
     processor_AB AB_4_2 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_2),
       .start_in   (start_in_4_2),
       .op_in      (op_in_4_2),
       .pivot_in   (pivot_in_4_2),
       .start_out  (start_out_4_2),
       .data_out   (data_out_4_2),
       .op_out     (op_out_4_2),
       .pivot_out  (pivot_out_4_2),
       .r          (r_4_2)
     );

  // row 4, col 3

     reg start_in_4_3;
     wire start_out_4_3;

     reg [1:0] op_in_4_3;
     wire [1:0] op_out_4_3;

     wire r_4_3;

     reg data_in_4_3;
     wire data_out_4_3;

     reg pivot_in_4_3;
     wire pivot_out_4_3;

     always @(posedge clk) begin
         op_in_4_3 <= op_out_4_2;
         pivot_in_4_3 <= pivot_out_4_2;
         start_in_4_3 <= start_out_4_2;
     end

     always @(posedge clk) begin
         data_in_4_3 <= data_out_3_3;
     end
  
     processor_AB AB_4_3 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_3),
       .start_in   (start_in_4_3),
       .op_in      (op_in_4_3),
       .pivot_in   (pivot_in_4_3),
       .start_out  (start_out_4_3),
       .data_out   (data_out_4_3),
       .op_out     (op_out_4_3),
       .pivot_out  (pivot_out_4_3),
       .r          (r_4_3)
     );

  // row 4, col 4

     reg start_in_4_4;
     wire start_out_4_4;

     reg [1:0] op_in_4_4;
     wire [1:0] op_out_4_4;

     wire r_4_4;

     reg data_in_4_4;
     wire data_out_4_4;

     reg pivot_in_4_4;
     wire pivot_out_4_4;

     always @(posedge clk) begin
         op_in_4_4 <= op_out_4_3;
         pivot_in_4_4 <= pivot_out_4_3;
         start_in_4_4 <= start_out_4_3;
     end

     always @(posedge clk) begin
         data_in_4_4 <= data_out_3_4;
     end
  
     processor_AB AB_4_4 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_4),
       .start_in   (start_in_4_4),
       .op_in      (op_in_4_4),
       .pivot_in   (pivot_in_4_4),
       .start_out  (start_out_4_4),
       .data_out   (data_out_4_4),
       .op_out     (op_out_4_4),
       .pivot_out  (pivot_out_4_4),
       .r          (r_4_4)
     );

  // row 4, col 5

     reg start_in_4_5;
     wire start_out_4_5;

     reg [1:0] op_in_4_5;
     wire [1:0] op_out_4_5;

     wire r_4_5;

     reg data_in_4_5;
     wire data_out_4_5;

     reg pivot_in_4_5;
     wire pivot_out_4_5;

     always @(posedge clk) begin
         op_in_4_5 <= op_out_4_4;
         pivot_in_4_5 <= pivot_out_4_4;
         start_in_4_5 <= start_out_4_4;
     end

     always @(posedge clk) begin
         data_in_4_5 <= data_out_3_5;
     end
  
     processor_AB AB_4_5 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_5),
       .start_in   (start_in_4_5),
       .op_in      (op_in_4_5),
       .pivot_in   (pivot_in_4_5),
       .start_out  (start_out_4_5),
       .data_out   (data_out_4_5),
       .op_out     (op_out_4_5),
       .pivot_out  (pivot_out_4_5),
       .r          (r_4_5)
     );

  // row 4, col 6

     reg start_in_4_6;
     wire start_out_4_6;

     reg [1:0] op_in_4_6;
     wire [1:0] op_out_4_6;

     wire r_4_6;

     reg data_in_4_6;
     wire data_out_4_6;

     reg pivot_in_4_6;
     wire pivot_out_4_6;

     always @(posedge clk) begin
         op_in_4_6 <= op_out_4_5;
         pivot_in_4_6 <= pivot_out_4_5;
         start_in_4_6 <= start_out_4_5;
     end

     always @(posedge clk) begin
         data_in_4_6 <= data_out_3_6;
     end
  
     processor_AB AB_4_6 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_6),
       .start_in   (start_in_4_6),
       .op_in      (op_in_4_6),
       .pivot_in   (pivot_in_4_6),
       .start_out  (start_out_4_6),
       .data_out   (data_out_4_6),
       .op_out     (op_out_4_6),
       .pivot_out  (pivot_out_4_6),
       .r          (r_4_6)
     );

  // row 4, col 7

     reg start_in_4_7;
     wire start_out_4_7;

     reg [1:0] op_in_4_7;
     wire [1:0] op_out_4_7;

     wire r_4_7;

     reg data_in_4_7;
     wire data_out_4_7;

     reg pivot_in_4_7;
     wire pivot_out_4_7;

     always @(posedge clk) begin
         op_in_4_7 <= op_out_4_6;
         pivot_in_4_7 <= pivot_out_4_6;
         start_in_4_7 <= start_out_4_6;
     end

     always @(posedge clk) begin
         data_in_4_7 <= data_out_3_7;
     end
  
     processor_AB AB_4_7 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_7),
       .start_in   (start_in_4_7),
       .op_in      (op_in_4_7),
       .pivot_in   (pivot_in_4_7),
       .start_out  (start_out_4_7),
       .data_out   (data_out_4_7),
       .op_out     (op_out_4_7),
       .pivot_out  (pivot_out_4_7),
       .r          (r_4_7)
     );

  // row 4, col 8

     reg start_in_4_8;
     wire start_out_4_8;

     reg [1:0] op_in_4_8;
     wire [1:0] op_out_4_8;

     wire r_4_8;

     reg data_in_4_8;
     wire data_out_4_8;

     reg pivot_in_4_8;
     wire pivot_out_4_8;

     always @(posedge clk) begin
         op_in_4_8 <= op_out_4_7;
         pivot_in_4_8 <= pivot_out_4_7;
         start_in_4_8 <= start_out_4_7;
     end

     always @(posedge clk) begin
         data_in_4_8 <= data_out_3_8;
     end
  
     processor_AB AB_4_8 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_8),
       .start_in   (start_in_4_8),
       .op_in      (op_in_4_8),
       .pivot_in   (pivot_in_4_8),
       .start_out  (start_out_4_8),
       .data_out   (data_out_4_8),
       .op_out     (op_out_4_8),
       .pivot_out  (pivot_out_4_8),
       .r          (r_4_8)
     );

  // row 4, col 9

     reg start_in_4_9;
     wire start_out_4_9;

     reg [1:0] op_in_4_9;
     wire [1:0] op_out_4_9;

     wire r_4_9;

     reg data_in_4_9;
     wire data_out_4_9;

     reg pivot_in_4_9;
     wire pivot_out_4_9;

     always @(posedge clk) begin
         op_in_4_9 <= op_out_4_8;
         pivot_in_4_9 <= pivot_out_4_8;
         start_in_4_9 <= start_out_4_8;
     end

     always @(posedge clk) begin
         data_in_4_9 <= data_out_3_9;
     end
  
     processor_AB AB_4_9 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_9),
       .start_in   (start_in_4_9),
       .op_in      (op_in_4_9),
       .pivot_in   (pivot_in_4_9),
       .start_out  (start_out_4_9),
       .data_out   (data_out_4_9),
       .op_out     (op_out_4_9),
       .pivot_out  (pivot_out_4_9),
       .r          (r_4_9)
     );

  // row 4, col 10

     reg start_in_4_10;
     wire start_out_4_10;

     reg [1:0] op_in_4_10;
     wire [1:0] op_out_4_10;

     wire r_4_10;

     reg data_in_4_10;
     wire data_out_4_10;

     reg pivot_in_4_10;
     wire pivot_out_4_10;

     always @(posedge clk) begin
         op_in_4_10 <= op_out_4_9;
         pivot_in_4_10 <= pivot_out_4_9;
         start_in_4_10 <= start_out_4_9;
     end

     always @(posedge clk) begin
         data_in_4_10 <= data_out_3_10;
     end
  
     processor_AB AB_4_10 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_10),
       .start_in   (start_in_4_10),
       .op_in      (op_in_4_10),
       .pivot_in   (pivot_in_4_10),
       .start_out  (start_out_4_10),
       .data_out   (data_out_4_10),
       .op_out     (op_out_4_10),
       .pivot_out  (pivot_out_4_10),
       .r          (r_4_10)
     );

  // row 4, col 11

     reg start_in_4_11;
     wire start_out_4_11;

     reg [1:0] op_in_4_11;
     wire [1:0] op_out_4_11;

     wire r_4_11;

     reg data_in_4_11;
     wire data_out_4_11;

     reg pivot_in_4_11;
     wire pivot_out_4_11;

     always @(posedge clk) begin
         op_in_4_11 <= op_out_4_10;
         pivot_in_4_11 <= pivot_out_4_10;
         start_in_4_11 <= start_out_4_10;
     end

     always @(posedge clk) begin
         data_in_4_11 <= data_out_3_11;
     end
  
     processor_AB AB_4_11 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_11),
       .start_in   (start_in_4_11),
       .op_in      (op_in_4_11),
       .pivot_in   (pivot_in_4_11),
       .start_out  (start_out_4_11),
       .data_out   (data_out_4_11),
       .op_out     (op_out_4_11),
       .pivot_out  (pivot_out_4_11),
       .r          (r_4_11)
     );

  // row 4, col 12

     reg start_in_4_12;
     wire start_out_4_12;

     reg [1:0] op_in_4_12;
     wire [1:0] op_out_4_12;

     wire r_4_12;

     reg data_in_4_12;
     wire data_out_4_12;

     reg pivot_in_4_12;
     wire pivot_out_4_12;

     always @(posedge clk) begin
         op_in_4_12 <= op_out_4_11;
         pivot_in_4_12 <= pivot_out_4_11;
         start_in_4_12 <= start_out_4_11;
     end

     always @(posedge clk) begin
         data_in_4_12 <= data_out_3_12;
     end
  
     processor_AB AB_4_12 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_12),
       .start_in   (start_in_4_12),
       .op_in      (op_in_4_12),
       .pivot_in   (pivot_in_4_12),
       .start_out  (start_out_4_12),
       .data_out   (data_out_4_12),
       .op_out     (op_out_4_12),
       .pivot_out  (pivot_out_4_12),
       .r          (r_4_12)
     );

  // row 4, col 13

     reg start_in_4_13;
     wire start_out_4_13;

     reg [1:0] op_in_4_13;
     wire [1:0] op_out_4_13;

     wire r_4_13;

     reg data_in_4_13;
     wire data_out_4_13;

     reg pivot_in_4_13;
     wire pivot_out_4_13;

     always @(posedge clk) begin
         op_in_4_13 <= op_out_4_12;
         pivot_in_4_13 <= pivot_out_4_12;
         start_in_4_13 <= start_out_4_12;
     end

     always @(posedge clk) begin
         data_in_4_13 <= data_out_3_13;
     end
  
     processor_AB AB_4_13 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_13),
       .start_in   (start_in_4_13),
       .op_in      (op_in_4_13),
       .pivot_in   (pivot_in_4_13),
       .start_out  (start_out_4_13),
       .data_out   (data_out_4_13),
       .op_out     (op_out_4_13),
       .pivot_out  (pivot_out_4_13),
       .r          (r_4_13)
     );

  // row 4, col 14

     reg start_in_4_14;
     wire start_out_4_14;

     reg [1:0] op_in_4_14;
     wire [1:0] op_out_4_14;

     wire r_4_14;

     reg data_in_4_14;
     wire data_out_4_14;

     reg pivot_in_4_14;
     wire pivot_out_4_14;

     always @(posedge clk) begin
         op_in_4_14 <= op_out_4_13;
         pivot_in_4_14 <= pivot_out_4_13;
         start_in_4_14 <= start_out_4_13;
     end

     always @(posedge clk) begin
         data_in_4_14 <= data_out_3_14;
     end
  
     processor_AB AB_4_14 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_14),
       .start_in   (start_in_4_14),
       .op_in      (op_in_4_14),
       .pivot_in   (pivot_in_4_14),
       .start_out  (start_out_4_14),
       .data_out   (data_out_4_14),
       .op_out     (op_out_4_14),
       .pivot_out  (pivot_out_4_14),
       .r          (r_4_14)
     );

  // row 4, col 15

     reg start_in_4_15;
     wire start_out_4_15;

     reg [1:0] op_in_4_15;
     wire [1:0] op_out_4_15;

     wire r_4_15;

     reg data_in_4_15;
     wire data_out_4_15;

     reg pivot_in_4_15;
     wire pivot_out_4_15;

     always @(posedge clk) begin
         op_in_4_15 <= op_out_4_14;
         pivot_in_4_15 <= pivot_out_4_14;
         start_in_4_15 <= start_out_4_14;
     end

     always @(posedge clk) begin
         data_in_4_15 <= data_out_3_15;
     end
  
     processor_AB AB_4_15 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_15),
       .start_in   (start_in_4_15),
       .op_in      (op_in_4_15),
       .pivot_in   (pivot_in_4_15),
       .start_out  (start_out_4_15),
       .data_out   (data_out_4_15),
       .op_out     (op_out_4_15),
       .pivot_out  (pivot_out_4_15),
       .r          (r_4_15)
     );

  // row 4, col 16

     reg start_in_4_16;
     wire start_out_4_16;

     reg [1:0] op_in_4_16;
     wire [1:0] op_out_4_16;

     wire r_4_16;

     reg data_in_4_16;
     wire data_out_4_16;

     reg pivot_in_4_16;
     wire pivot_out_4_16;

     always @(posedge clk) begin
         op_in_4_16 <= op_out_4_15;
         pivot_in_4_16 <= pivot_out_4_15;
         start_in_4_16 <= start_out_4_15;
     end

     always @(posedge clk) begin
         data_in_4_16 <= data_out_3_16;
     end
  
     processor_AB AB_4_16 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_16),
       .start_in   (start_in_4_16),
       .op_in      (op_in_4_16),
       .pivot_in   (pivot_in_4_16),
       .start_out  (start_out_4_16),
       .data_out   (data_out_4_16),
       .op_out     (op_out_4_16),
       .pivot_out  (pivot_out_4_16),
       .r          (r_4_16)
     );

  // row 4, col 17

     reg start_in_4_17;
     wire start_out_4_17;

     reg [1:0] op_in_4_17;
     wire [1:0] op_out_4_17;

     wire r_4_17;

     reg data_in_4_17;
     wire data_out_4_17;

     reg pivot_in_4_17;
     wire pivot_out_4_17;

     always @(posedge clk) begin
         op_in_4_17 <= op_out_4_16;
         pivot_in_4_17 <= pivot_out_4_16;
         start_in_4_17 <= start_out_4_16;
     end

     always @(posedge clk) begin
         data_in_4_17 <= data_out_3_17;
     end
  
     processor_AB AB_4_17 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_17),
       .start_in   (start_in_4_17),
       .op_in      (op_in_4_17),
       .pivot_in   (pivot_in_4_17),
       .start_out  (start_out_4_17),
       .data_out   (data_out_4_17),
       .op_out     (op_out_4_17),
       .pivot_out  (pivot_out_4_17),
       .r          (r_4_17)
     );

  // row 4, col 18

     reg start_in_4_18;
     wire start_out_4_18;

     reg [1:0] op_in_4_18;
     wire [1:0] op_out_4_18;

     wire r_4_18;

     reg data_in_4_18;
     wire data_out_4_18;

     reg pivot_in_4_18;
     wire pivot_out_4_18;

     always @(posedge clk) begin
         op_in_4_18 <= op_out_4_17;
         pivot_in_4_18 <= pivot_out_4_17;
         start_in_4_18 <= start_out_4_17;
     end

     always @(posedge clk) begin
         data_in_4_18 <= data_out_3_18;
     end
  
     processor_AB AB_4_18 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_18),
       .start_in   (start_in_4_18),
       .op_in      (op_in_4_18),
       .pivot_in   (pivot_in_4_18),
       .start_out  (start_out_4_18),
       .data_out   (data_out_4_18),
       .op_out     (op_out_4_18),
       .pivot_out  (pivot_out_4_18),
       .r          (r_4_18)
     );

  // row 4, col 19

     reg start_in_4_19;
     wire start_out_4_19;

     reg [1:0] op_in_4_19;
     wire [1:0] op_out_4_19;

     wire r_4_19;

     reg data_in_4_19;
     wire data_out_4_19;

     reg pivot_in_4_19;
     wire pivot_out_4_19;

     always @(posedge clk) begin
         op_in_4_19 <= op_out_4_18;
         pivot_in_4_19 <= pivot_out_4_18;
         start_in_4_19 <= start_out_4_18;
     end

     always @(posedge clk) begin
         data_in_4_19 <= data_out_3_19;
     end
  
     processor_AB AB_4_19 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_19),
       .start_in   (start_in_4_19),
       .op_in      (op_in_4_19),
       .pivot_in   (pivot_in_4_19),
       .start_out  (start_out_4_19),
       .data_out   (data_out_4_19),
       .op_out     (op_out_4_19),
       .pivot_out  (pivot_out_4_19),
       .r          (r_4_19)
     );

  // row 4, col 20

     reg start_in_4_20;
     wire start_out_4_20;

     reg [1:0] op_in_4_20;
     wire [1:0] op_out_4_20;

     wire r_4_20;

     reg data_in_4_20;
     wire data_out_4_20;

     reg pivot_in_4_20;
     wire pivot_out_4_20;

     always @(posedge clk) begin
         op_in_4_20 <= op_out_4_19;
         pivot_in_4_20 <= pivot_out_4_19;
         start_in_4_20 <= start_out_4_19;
     end

     always @(posedge clk) begin
         data_in_4_20 <= data_out_3_20;
     end
  
     processor_AB AB_4_20 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_20),
       .start_in   (start_in_4_20),
       .op_in      (op_in_4_20),
       .pivot_in   (pivot_in_4_20),
       .start_out  (start_out_4_20),
       .data_out   (data_out_4_20),
       .op_out     (op_out_4_20),
       .pivot_out  (pivot_out_4_20),
       .r          (r_4_20)
     );

  // row 4, col 21

     reg start_in_4_21;
     wire start_out_4_21;

     reg [1:0] op_in_4_21;
     wire [1:0] op_out_4_21;

     wire r_4_21;

     reg data_in_4_21;
     wire data_out_4_21;

     reg pivot_in_4_21;
     wire pivot_out_4_21;

     always @(posedge clk) begin
         op_in_4_21 <= op_out_4_20;
         pivot_in_4_21 <= pivot_out_4_20;
         start_in_4_21 <= start_out_4_20;
     end

     always @(posedge clk) begin
         data_in_4_21 <= data_out_3_21;
     end
  
     processor_AB AB_4_21 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_21),
       .start_in   (start_in_4_21),
       .op_in      (op_in_4_21),
       .pivot_in   (pivot_in_4_21),
       .start_out  (start_out_4_21),
       .data_out   (data_out_4_21),
       .op_out     (op_out_4_21),
       .pivot_out  (pivot_out_4_21),
       .r          (r_4_21)
     );

  // row 4, col 22

     reg start_in_4_22;
     wire start_out_4_22;

     reg [1:0] op_in_4_22;
     wire [1:0] op_out_4_22;

     wire r_4_22;

     reg data_in_4_22;
     wire data_out_4_22;

     reg pivot_in_4_22;
     wire pivot_out_4_22;

     always @(posedge clk) begin
         op_in_4_22 <= op_out_4_21;
         pivot_in_4_22 <= pivot_out_4_21;
         start_in_4_22 <= start_out_4_21;
     end

     always @(posedge clk) begin
         data_in_4_22 <= data_out_3_22;
     end
  
     processor_AB AB_4_22 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_22),
       .start_in   (start_in_4_22),
       .op_in      (op_in_4_22),
       .pivot_in   (pivot_in_4_22),
       .start_out  (start_out_4_22),
       .data_out   (data_out_4_22),
       .op_out     (op_out_4_22),
       .pivot_out  (pivot_out_4_22),
       .r          (r_4_22)
     );

  // row 4, col 23

     reg start_in_4_23;
     wire start_out_4_23;

     reg [1:0] op_in_4_23;
     wire [1:0] op_out_4_23;

     wire r_4_23;

     reg data_in_4_23;
     wire data_out_4_23;

     reg pivot_in_4_23;
     wire pivot_out_4_23;

     always @(posedge clk) begin
         op_in_4_23 <= op_out_4_22;
         pivot_in_4_23 <= pivot_out_4_22;
         start_in_4_23 <= start_out_4_22;
     end

     always @(posedge clk) begin
         data_in_4_23 <= data_out_3_23;
     end
  
     processor_AB AB_4_23 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_23),
       .start_in   (start_in_4_23),
       .op_in      (op_in_4_23),
       .pivot_in   (pivot_in_4_23),
       .start_out  (start_out_4_23),
       .data_out   (data_out_4_23),
       .op_out     (op_out_4_23),
       .pivot_out  (pivot_out_4_23),
       .r          (r_4_23)
     );

  // row 4, col 24

     reg start_in_4_24;
     wire start_out_4_24;

     reg [1:0] op_in_4_24;
     wire [1:0] op_out_4_24;

     wire r_4_24;

     reg data_in_4_24;
     wire data_out_4_24;

     reg pivot_in_4_24;
     wire pivot_out_4_24;

     always @(posedge clk) begin
         op_in_4_24 <= op_out_4_23;
         pivot_in_4_24 <= pivot_out_4_23;
         start_in_4_24 <= start_out_4_23;
     end

     always @(posedge clk) begin
         data_in_4_24 <= data_out_3_24;
     end
  
     processor_AB AB_4_24 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_24),
       .start_in   (start_in_4_24),
       .op_in      (op_in_4_24),
       .pivot_in   (pivot_in_4_24),
       .start_out  (start_out_4_24),
       .data_out   (data_out_4_24),
       .op_out     (op_out_4_24),
       .pivot_out  (pivot_out_4_24),
       .r          (r_4_24)
     );

  // row 4, col 25

     reg start_in_4_25;
     wire start_out_4_25;

     reg [1:0] op_in_4_25;
     wire [1:0] op_out_4_25;

     wire r_4_25;

     reg data_in_4_25;
     wire data_out_4_25;

     reg pivot_in_4_25;
     wire pivot_out_4_25;

     always @(posedge clk) begin
         op_in_4_25 <= op_out_4_24;
         pivot_in_4_25 <= pivot_out_4_24;
         start_in_4_25 <= start_out_4_24;
     end

     always @(posedge clk) begin
         data_in_4_25 <= data_out_3_25;
     end
  
     processor_AB AB_4_25 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_25),
       .start_in   (start_in_4_25),
       .op_in      (op_in_4_25),
       .pivot_in   (pivot_in_4_25),
       .start_out  (start_out_4_25),
       .data_out   (data_out_4_25),
       .op_out     (op_out_4_25),
       .pivot_out  (pivot_out_4_25),
       .r          (r_4_25)
     );

  // row 4, col 26

     reg start_in_4_26;
     wire start_out_4_26;

     reg [1:0] op_in_4_26;
     wire [1:0] op_out_4_26;

     wire r_4_26;

     reg data_in_4_26;
     wire data_out_4_26;

     reg pivot_in_4_26;
     wire pivot_out_4_26;

     always @(posedge clk) begin
         op_in_4_26 <= op_out_4_25;
         pivot_in_4_26 <= pivot_out_4_25;
         start_in_4_26 <= start_out_4_25;
     end

     always @(posedge clk) begin
         data_in_4_26 <= data_out_3_26;
     end
  
     processor_AB AB_4_26 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_26),
       .start_in   (start_in_4_26),
       .op_in      (op_in_4_26),
       .pivot_in   (pivot_in_4_26),
       .start_out  (start_out_4_26),
       .data_out   (data_out_4_26),
       .op_out     (op_out_4_26),
       .pivot_out  (pivot_out_4_26),
       .r          (r_4_26)
     );

  // row 4, col 27

     reg start_in_4_27;
     wire start_out_4_27;

     reg [1:0] op_in_4_27;
     wire [1:0] op_out_4_27;

     wire r_4_27;

     reg data_in_4_27;
     wire data_out_4_27;

     reg pivot_in_4_27;
     wire pivot_out_4_27;

     always @(posedge clk) begin
         op_in_4_27 <= op_out_4_26;
         pivot_in_4_27 <= pivot_out_4_26;
         start_in_4_27 <= start_out_4_26;
     end

     always @(posedge clk) begin
         data_in_4_27 <= data_out_3_27;
     end
  
     processor_AB AB_4_27 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_27),
       .start_in   (start_in_4_27),
       .op_in      (op_in_4_27),
       .pivot_in   (pivot_in_4_27),
       .start_out  (start_out_4_27),
       .data_out   (data_out_4_27),
       .op_out     (op_out_4_27),
       .pivot_out  (pivot_out_4_27),
       .r          (r_4_27)
     );

  // row 4, col 28

     reg start_in_4_28;
     wire start_out_4_28;

     reg [1:0] op_in_4_28;
     wire [1:0] op_out_4_28;

     wire r_4_28;

     reg data_in_4_28;
     wire data_out_4_28;

     reg pivot_in_4_28;
     wire pivot_out_4_28;

     always @(posedge clk) begin
         op_in_4_28 <= op_out_4_27;
         pivot_in_4_28 <= pivot_out_4_27;
         start_in_4_28 <= start_out_4_27;
     end

     always @(posedge clk) begin
         data_in_4_28 <= data_out_3_28;
     end
  
     processor_AB AB_4_28 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_28),
       .start_in   (start_in_4_28),
       .op_in      (op_in_4_28),
       .pivot_in   (pivot_in_4_28),
       .start_out  (start_out_4_28),
       .data_out   (data_out_4_28),
       .op_out     (op_out_4_28),
       .pivot_out  (pivot_out_4_28),
       .r          (r_4_28)
     );

  // row 4, col 29

     reg start_in_4_29;
     wire start_out_4_29;

     reg [1:0] op_in_4_29;
     wire [1:0] op_out_4_29;

     wire r_4_29;

     reg data_in_4_29;
     wire data_out_4_29;

     reg pivot_in_4_29;
     wire pivot_out_4_29;

     always @(posedge clk) begin
         op_in_4_29 <= op_out_4_28;
         pivot_in_4_29 <= pivot_out_4_28;
         start_in_4_29 <= start_out_4_28;
     end

     always @(posedge clk) begin
         data_in_4_29 <= data_out_3_29;
     end
  
     processor_AB AB_4_29 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_29),
       .start_in   (start_in_4_29),
       .op_in      (op_in_4_29),
       .pivot_in   (pivot_in_4_29),
       .start_out  (start_out_4_29),
       .data_out   (data_out_4_29),
       .op_out     (op_out_4_29),
       .pivot_out  (pivot_out_4_29),
       .r          (r_4_29)
     );

  // row 4, col 30

     reg start_in_4_30;
     wire start_out_4_30;

     reg [1:0] op_in_4_30;
     wire [1:0] op_out_4_30;

     wire r_4_30;

     reg data_in_4_30;
     wire data_out_4_30;

     reg pivot_in_4_30;
     wire pivot_out_4_30;

     always @(posedge clk) begin
         op_in_4_30 <= op_out_4_29;
         pivot_in_4_30 <= pivot_out_4_29;
         start_in_4_30 <= start_out_4_29;
     end

     always @(posedge clk) begin
         data_in_4_30 <= data_out_3_30;
     end
  
     processor_AB AB_4_30 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_30),
       .start_in   (start_in_4_30),
       .op_in      (op_in_4_30),
       .pivot_in   (pivot_in_4_30),
       .start_out  (start_out_4_30),
       .data_out   (data_out_4_30),
       .op_out     (op_out_4_30),
       .pivot_out  (pivot_out_4_30),
       .r          (r_4_30)
     );

  // row 4, col 31

     reg start_in_4_31;
     wire start_out_4_31;

     reg [1:0] op_in_4_31;
     wire [1:0] op_out_4_31;

     wire r_4_31;

     reg data_in_4_31;
     wire data_out_4_31;

     reg pivot_in_4_31;
     wire pivot_out_4_31;

     always @(posedge clk) begin
         op_in_4_31 <= op_out_4_30;
         pivot_in_4_31 <= pivot_out_4_30;
         start_in_4_31 <= start_out_4_30;
     end

     always @(posedge clk) begin
         data_in_4_31 <= data_out_3_31;
     end
  
     processor_AB AB_4_31 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_31),
       .start_in   (start_in_4_31),
       .op_in      (op_in_4_31),
       .pivot_in   (pivot_in_4_31),
       .start_out  (start_out_4_31),
       .data_out   (data_out_4_31),
       .op_out     (op_out_4_31),
       .pivot_out  (pivot_out_4_31),
       .r          (r_4_31)
     );

  // row 4, col 32

     reg start_in_4_32;
     wire start_out_4_32;

     reg [1:0] op_in_4_32;
     wire [1:0] op_out_4_32;

     wire r_4_32;

     reg data_in_4_32;
     wire data_out_4_32;

     reg pivot_in_4_32;
     wire pivot_out_4_32;

     always @(posedge clk) begin
         op_in_4_32 <= op_out_4_31;
         pivot_in_4_32 <= pivot_out_4_31;
         start_in_4_32 <= start_out_4_31;
     end

     always @(posedge clk) begin
         data_in_4_32 <= data_out_3_32;
     end
  
     processor_AB AB_4_32 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_32),
       .start_in   (start_in_4_32),
       .op_in      (op_in_4_32),
       .pivot_in   (pivot_in_4_32),
       .start_out  (start_out_4_32),
       .data_out   (data_out_4_32),
       .op_out     (op_out_4_32),
       .pivot_out  (pivot_out_4_32),
       .r          (r_4_32)
     );

  // row 4, col 33

     reg start_in_4_33;
     wire start_out_4_33;

     reg [1:0] op_in_4_33;
     wire [1:0] op_out_4_33;

     wire r_4_33;

     reg data_in_4_33;
     wire data_out_4_33;

     reg pivot_in_4_33;
     wire pivot_out_4_33;

     always @(posedge clk) begin
         op_in_4_33 <= op_out_4_32;
         pivot_in_4_33 <= pivot_out_4_32;
         start_in_4_33 <= start_out_4_32;
     end

     always @(posedge clk) begin
         data_in_4_33 <= data_out_3_33;
     end
  
     processor_AB AB_4_33 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_33),
       .start_in   (start_in_4_33),
       .op_in      (op_in_4_33),
       .pivot_in   (pivot_in_4_33),
       .start_out  (start_out_4_33),
       .data_out   (data_out_4_33),
       .op_out     (op_out_4_33),
       .pivot_out  (pivot_out_4_33),
       .r          (r_4_33)
     );

  // row 4, col 34

     reg start_in_4_34;
     wire start_out_4_34;

     reg [1:0] op_in_4_34;
     wire [1:0] op_out_4_34;

     wire r_4_34;

     reg data_in_4_34;
     wire data_out_4_34;

     reg pivot_in_4_34;
     wire pivot_out_4_34;

     always @(posedge clk) begin
         op_in_4_34 <= op_out_4_33;
         pivot_in_4_34 <= pivot_out_4_33;
         start_in_4_34 <= start_out_4_33;
     end

     always @(posedge clk) begin
         data_in_4_34 <= data_out_3_34;
     end
  
     processor_AB AB_4_34 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_34),
       .start_in   (start_in_4_34),
       .op_in      (op_in_4_34),
       .pivot_in   (pivot_in_4_34),
       .start_out  (start_out_4_34),
       .data_out   (data_out_4_34),
       .op_out     (op_out_4_34),
       .pivot_out  (pivot_out_4_34),
       .r          (r_4_34)
     );

  // row 4, col 35

     reg start_in_4_35;
     wire start_out_4_35;

     reg [1:0] op_in_4_35;
     wire [1:0] op_out_4_35;

     wire r_4_35;

     reg data_in_4_35;
     wire data_out_4_35;

     reg pivot_in_4_35;
     wire pivot_out_4_35;

     always @(posedge clk) begin
         op_in_4_35 <= op_out_4_34;
         pivot_in_4_35 <= pivot_out_4_34;
         start_in_4_35 <= start_out_4_34;
     end

     always @(posedge clk) begin
         data_in_4_35 <= data_out_3_35;
     end
  
     processor_AB AB_4_35 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_35),
       .start_in   (start_in_4_35),
       .op_in      (op_in_4_35),
       .pivot_in   (pivot_in_4_35),
       .start_out  (start_out_4_35),
       .data_out   (data_out_4_35),
       .op_out     (op_out_4_35),
       .pivot_out  (pivot_out_4_35),
       .r          (r_4_35)
     );

  // row 4, col 36

     reg start_in_4_36;
     wire start_out_4_36;

     reg [1:0] op_in_4_36;
     wire [1:0] op_out_4_36;

     wire r_4_36;

     reg data_in_4_36;
     wire data_out_4_36;

     reg pivot_in_4_36;
     wire pivot_out_4_36;

     always @(posedge clk) begin
         op_in_4_36 <= op_out_4_35;
         pivot_in_4_36 <= pivot_out_4_35;
         start_in_4_36 <= start_out_4_35;
     end

     always @(posedge clk) begin
         data_in_4_36 <= data_out_3_36;
     end
  
     processor_AB AB_4_36 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_36),
       .start_in   (start_in_4_36),
       .op_in      (op_in_4_36),
       .pivot_in   (pivot_in_4_36),
       .start_out  (start_out_4_36),
       .data_out   (data_out_4_36),
       .op_out     (op_out_4_36),
       .pivot_out  (pivot_out_4_36),
       .r          (r_4_36)
     );

  // row 4, col 37

     reg start_in_4_37;
     wire start_out_4_37;

     reg [1:0] op_in_4_37;
     wire [1:0] op_out_4_37;

     wire r_4_37;

     reg data_in_4_37;
     wire data_out_4_37;

     reg pivot_in_4_37;
     wire pivot_out_4_37;

     always @(posedge clk) begin
         op_in_4_37 <= op_out_4_36;
         pivot_in_4_37 <= pivot_out_4_36;
         start_in_4_37 <= start_out_4_36;
     end

     always @(posedge clk) begin
         data_in_4_37 <= data_out_3_37;
     end
  
     processor_AB AB_4_37 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_37),
       .start_in   (start_in_4_37),
       .op_in      (op_in_4_37),
       .pivot_in   (pivot_in_4_37),
       .start_out  (start_out_4_37),
       .data_out   (data_out_4_37),
       .op_out     (op_out_4_37),
       .pivot_out  (pivot_out_4_37),
       .r          (r_4_37)
     );

  // row 4, col 38

     reg start_in_4_38;
     wire start_out_4_38;

     reg [1:0] op_in_4_38;
     wire [1:0] op_out_4_38;

     wire r_4_38;

     reg data_in_4_38;
     wire data_out_4_38;

     reg pivot_in_4_38;
     wire pivot_out_4_38;

     always @(posedge clk) begin
         op_in_4_38 <= op_out_4_37;
         pivot_in_4_38 <= pivot_out_4_37;
         start_in_4_38 <= start_out_4_37;
     end

     always @(posedge clk) begin
         data_in_4_38 <= data_out_3_38;
     end
  
     processor_AB AB_4_38 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_38),
       .start_in   (start_in_4_38),
       .op_in      (op_in_4_38),
       .pivot_in   (pivot_in_4_38),
       .start_out  (start_out_4_38),
       .data_out   (data_out_4_38),
       .op_out     (op_out_4_38),
       .pivot_out  (pivot_out_4_38),
       .r          (r_4_38)
     );

  // row 4, col 39

     reg start_in_4_39;
     wire start_out_4_39;

     reg [1:0] op_in_4_39;
     wire [1:0] op_out_4_39;

     wire r_4_39;

     reg data_in_4_39;
     wire data_out_4_39;

     reg pivot_in_4_39;
     wire pivot_out_4_39;

     always @(posedge clk) begin
         op_in_4_39 <= op_out_4_38;
         pivot_in_4_39 <= pivot_out_4_38;
         start_in_4_39 <= start_out_4_38;
     end

     always @(posedge clk) begin
         data_in_4_39 <= data_out_3_39;
     end
  
     processor_AB AB_4_39 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_39),
       .start_in   (start_in_4_39),
       .op_in      (op_in_4_39),
       .pivot_in   (pivot_in_4_39),
       .start_out  (start_out_4_39),
       .data_out   (data_out_4_39),
       .op_out     (op_out_4_39),
       .pivot_out  (pivot_out_4_39),
       .r          (r_4_39)
     );

  // row 4, col 40

     reg start_in_4_40;
     wire start_out_4_40;

     reg [1:0] op_in_4_40;
     wire [1:0] op_out_4_40;

     wire r_4_40;

     reg data_in_4_40;
     wire data_out_4_40;

     reg pivot_in_4_40;
     wire pivot_out_4_40;

     always @(posedge clk) begin
         op_in_4_40 <= op_out_4_39;
         pivot_in_4_40 <= pivot_out_4_39;
         start_in_4_40 <= start_out_4_39;
     end

     always @(posedge clk) begin
         data_in_4_40 <= data_out_3_40;
     end
  
     processor_AB AB_4_40 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_40),
       .start_in   (start_in_4_40),
       .op_in      (op_in_4_40),
       .pivot_in   (pivot_in_4_40),
       .start_out  (start_out_4_40),
       .data_out   (data_out_4_40),
       .op_out     (op_out_4_40),
       .pivot_out  (pivot_out_4_40),
       .r          (r_4_40)
     );

  // row 4, col 41

     reg start_in_4_41;
     wire start_out_4_41;

     reg [1:0] op_in_4_41;
     wire [1:0] op_out_4_41;

     wire r_4_41;

     reg data_in_4_41;
     wire data_out_4_41;

     reg pivot_in_4_41;
     wire pivot_out_4_41;

     always @(posedge clk) begin
         op_in_4_41 <= op_out_4_40;
         pivot_in_4_41 <= pivot_out_4_40;
         start_in_4_41 <= start_out_4_40;
     end

     always @(posedge clk) begin
         data_in_4_41 <= data_out_3_41;
     end
  
     processor_AB AB_4_41 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_41),
       .start_in   (start_in_4_41),
       .op_in      (op_in_4_41),
       .pivot_in   (pivot_in_4_41),
       .start_out  (start_out_4_41),
       .data_out   (data_out_4_41),
       .op_out     (op_out_4_41),
       .pivot_out  (pivot_out_4_41),
       .r          (r_4_41)
     );

  // row 4, col 42

     reg start_in_4_42;
     wire start_out_4_42;

     reg [1:0] op_in_4_42;
     wire [1:0] op_out_4_42;

     wire r_4_42;

     reg data_in_4_42;
     wire data_out_4_42;

     reg pivot_in_4_42;
     wire pivot_out_4_42;

     always @(posedge clk) begin
         op_in_4_42 <= op_out_4_41;
         pivot_in_4_42 <= pivot_out_4_41;
         start_in_4_42 <= start_out_4_41;
     end

     always @(posedge clk) begin
         data_in_4_42 <= data_out_3_42;
     end
  
     processor_AB AB_4_42 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_42),
       .start_in   (start_in_4_42),
       .op_in      (op_in_4_42),
       .pivot_in   (pivot_in_4_42),
       .start_out  (start_out_4_42),
       .data_out   (data_out_4_42),
       .op_out     (op_out_4_42),
       .pivot_out  (pivot_out_4_42),
       .r          (r_4_42)
     );

  // row 4, col 43

     reg start_in_4_43;
     wire start_out_4_43;

     reg [1:0] op_in_4_43;
     wire [1:0] op_out_4_43;

     wire r_4_43;

     reg data_in_4_43;
     wire data_out_4_43;

     reg pivot_in_4_43;
     wire pivot_out_4_43;

     always @(posedge clk) begin
         op_in_4_43 <= op_out_4_42;
         pivot_in_4_43 <= pivot_out_4_42;
         start_in_4_43 <= start_out_4_42;
     end

     always @(posedge clk) begin
         data_in_4_43 <= data_out_3_43;
     end
  
     processor_AB AB_4_43 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_43),
       .start_in   (start_in_4_43),
       .op_in      (op_in_4_43),
       .pivot_in   (pivot_in_4_43),
       .start_out  (start_out_4_43),
       .data_out   (data_out_4_43),
       .op_out     (op_out_4_43),
       .pivot_out  (pivot_out_4_43),
       .r          (r_4_43)
     );

  // row 4, col 44

     reg start_in_4_44;
     wire start_out_4_44;

     reg [1:0] op_in_4_44;
     wire [1:0] op_out_4_44;

     wire r_4_44;

     reg data_in_4_44;
     wire data_out_4_44;

     reg pivot_in_4_44;
     wire pivot_out_4_44;

     always @(posedge clk) begin
         op_in_4_44 <= op_out_4_43;
         pivot_in_4_44 <= pivot_out_4_43;
         start_in_4_44 <= start_out_4_43;
     end

     always @(posedge clk) begin
         data_in_4_44 <= data_out_3_44;
     end
  
     processor_AB AB_4_44 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_44),
       .start_in   (start_in_4_44),
       .op_in      (op_in_4_44),
       .pivot_in   (pivot_in_4_44),
       .start_out  (start_out_4_44),
       .data_out   (data_out_4_44),
       .op_out     (op_out_4_44),
       .pivot_out  (pivot_out_4_44),
       .r          (r_4_44)
     );

  // row 4, col 45

     reg start_in_4_45;
     wire start_out_4_45;

     reg [1:0] op_in_4_45;
     wire [1:0] op_out_4_45;

     wire r_4_45;

     reg data_in_4_45;
     wire data_out_4_45;

     reg pivot_in_4_45;
     wire pivot_out_4_45;

     always @(posedge clk) begin
         op_in_4_45 <= op_out_4_44;
         pivot_in_4_45 <= pivot_out_4_44;
         start_in_4_45 <= start_out_4_44;
     end

     always @(posedge clk) begin
         data_in_4_45 <= data_out_3_45;
     end
  
     processor_AB AB_4_45 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_45),
       .start_in   (start_in_4_45),
       .op_in      (op_in_4_45),
       .pivot_in   (pivot_in_4_45),
       .start_out  (start_out_4_45),
       .data_out   (data_out_4_45),
       .op_out     (op_out_4_45),
       .pivot_out  (pivot_out_4_45),
       .r          (r_4_45)
     );

  // row 4, col 46

     reg start_in_4_46;
     wire start_out_4_46;

     reg [1:0] op_in_4_46;
     wire [1:0] op_out_4_46;

     wire r_4_46;

     reg data_in_4_46;
     wire data_out_4_46;

     reg pivot_in_4_46;
     wire pivot_out_4_46;

     always @(posedge clk) begin
         op_in_4_46 <= op_out_4_45;
         pivot_in_4_46 <= pivot_out_4_45;
         start_in_4_46 <= start_out_4_45;
     end

     always @(posedge clk) begin
         data_in_4_46 <= data_out_3_46;
     end
  
     processor_AB AB_4_46 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_46),
       .start_in   (start_in_4_46),
       .op_in      (op_in_4_46),
       .pivot_in   (pivot_in_4_46),
       .start_out  (start_out_4_46),
       .data_out   (data_out_4_46),
       .op_out     (op_out_4_46),
       .pivot_out  (pivot_out_4_46),
       .r          (r_4_46)
     );

  // row 4, col 47

     reg start_in_4_47;
     wire start_out_4_47;

     reg [1:0] op_in_4_47;
     wire [1:0] op_out_4_47;

     wire r_4_47;

     reg data_in_4_47;
     wire data_out_4_47;

     reg pivot_in_4_47;
     wire pivot_out_4_47;

     always @(posedge clk) begin
         op_in_4_47 <= op_out_4_46;
         pivot_in_4_47 <= pivot_out_4_46;
         start_in_4_47 <= start_out_4_46;
     end

     always @(posedge clk) begin
         data_in_4_47 <= data_out_3_47;
     end
  
     processor_AB AB_4_47 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_47),
       .start_in   (start_in_4_47),
       .op_in      (op_in_4_47),
       .pivot_in   (pivot_in_4_47),
       .start_out  (start_out_4_47),
       .data_out   (data_out_4_47),
       .op_out     (op_out_4_47),
       .pivot_out  (pivot_out_4_47),
       .r          (r_4_47)
     );

  // row 4, col 48

     reg start_in_4_48;
     wire start_out_4_48;

     reg [1:0] op_in_4_48;
     wire [1:0] op_out_4_48;

     wire r_4_48;

     reg data_in_4_48;
     wire data_out_4_48;

     reg pivot_in_4_48;
     wire pivot_out_4_48;

     always @(posedge clk) begin
         op_in_4_48 <= op_out_4_47;
         pivot_in_4_48 <= pivot_out_4_47;
         start_in_4_48 <= start_out_4_47;
     end

     always @(posedge clk) begin
         data_in_4_48 <= data_out_3_48;
     end
  
     processor_AB AB_4_48 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_48),
       .start_in   (start_in_4_48),
       .op_in      (op_in_4_48),
       .pivot_in   (pivot_in_4_48),
       .start_out  (start_out_4_48),
       .data_out   (data_out_4_48),
       .op_out     (op_out_4_48),
       .pivot_out  (pivot_out_4_48),
       .r          (r_4_48)
     );

  // row 4, col 49

     reg start_in_4_49;
     wire start_out_4_49;

     reg [1:0] op_in_4_49;
     wire [1:0] op_out_4_49;

     wire r_4_49;

     reg data_in_4_49;
     wire data_out_4_49;

     reg pivot_in_4_49;
     wire pivot_out_4_49;

     always @(posedge clk) begin
         op_in_4_49 <= op_out_4_48;
         pivot_in_4_49 <= pivot_out_4_48;
         start_in_4_49 <= start_out_4_48;
     end

     always @(posedge clk) begin
         data_in_4_49 <= data_out_3_49;
     end
  
     processor_AB AB_4_49 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_49),
       .start_in   (start_in_4_49),
       .op_in      (op_in_4_49),
       .pivot_in   (pivot_in_4_49),
       .start_out  (start_out_4_49),
       .data_out   (data_out_4_49),
       .op_out     (op_out_4_49),
       .pivot_out  (pivot_out_4_49),
       .r          (r_4_49)
     );

  // row 4, col 50

     reg start_in_4_50;
     wire start_out_4_50;

     reg [1:0] op_in_4_50;
     wire [1:0] op_out_4_50;

     wire r_4_50;

     reg data_in_4_50;
     wire data_out_4_50;

     reg pivot_in_4_50;
     wire pivot_out_4_50;

     always @(posedge clk) begin
         op_in_4_50 <= op_out_4_49;
         pivot_in_4_50 <= pivot_out_4_49;
         start_in_4_50 <= start_out_4_49;
     end

     always @(posedge clk) begin
         data_in_4_50 <= data_out_3_50;
     end
  
     processor_AB AB_4_50 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_50),
       .start_in   (start_in_4_50),
       .op_in      (op_in_4_50),
       .pivot_in   (pivot_in_4_50),
       .start_out  (start_out_4_50),
       .data_out   (data_out_4_50),
       .op_out     (op_out_4_50),
       .pivot_out  (pivot_out_4_50),
       .r          (r_4_50)
     );

  // row 4, col 51

     reg start_in_4_51;
     wire start_out_4_51;

     reg [1:0] op_in_4_51;
     wire [1:0] op_out_4_51;

     wire r_4_51;

     reg data_in_4_51;
     wire data_out_4_51;

     reg pivot_in_4_51;
     wire pivot_out_4_51;

     always @(posedge clk) begin
         op_in_4_51 <= op_out_4_50;
         pivot_in_4_51 <= pivot_out_4_50;
         start_in_4_51 <= start_out_4_50;
     end

     always @(posedge clk) begin
         data_in_4_51 <= data_out_3_51;
     end
  
     processor_AB AB_4_51 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_51),
       .start_in   (start_in_4_51),
       .op_in      (op_in_4_51),
       .pivot_in   (pivot_in_4_51),
       .start_out  (start_out_4_51),
       .data_out   (data_out_4_51),
       .op_out     (op_out_4_51),
       .pivot_out  (pivot_out_4_51),
       .r          (r_4_51)
     );

  // row 4, col 52

     reg start_in_4_52;
     wire start_out_4_52;

     reg [1:0] op_in_4_52;
     wire [1:0] op_out_4_52;

     wire r_4_52;

     reg data_in_4_52;
     wire data_out_4_52;

     reg pivot_in_4_52;
     wire pivot_out_4_52;

     always @(posedge clk) begin
         op_in_4_52 <= op_out_4_51;
         pivot_in_4_52 <= pivot_out_4_51;
         start_in_4_52 <= start_out_4_51;
     end

     always @(posedge clk) begin
         data_in_4_52 <= data_out_3_52;
     end
  
     processor_AB AB_4_52 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_52),
       .start_in   (start_in_4_52),
       .op_in      (op_in_4_52),
       .pivot_in   (pivot_in_4_52),
       .start_out  (start_out_4_52),
       .data_out   (data_out_4_52),
       .op_out     (op_out_4_52),
       .pivot_out  (pivot_out_4_52),
       .r          (r_4_52)
     );

  // row 4, col 53

     reg start_in_4_53;
     wire start_out_4_53;

     reg [1:0] op_in_4_53;
     wire [1:0] op_out_4_53;

     wire r_4_53;

     reg data_in_4_53;
     wire data_out_4_53;

     reg pivot_in_4_53;
     wire pivot_out_4_53;

     always @(posedge clk) begin
         op_in_4_53 <= op_out_4_52;
         pivot_in_4_53 <= pivot_out_4_52;
         start_in_4_53 <= start_out_4_52;
     end

     always @(posedge clk) begin
         data_in_4_53 <= data_out_3_53;
     end
  
     processor_AB AB_4_53 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_53),
       .start_in   (start_in_4_53),
       .op_in      (op_in_4_53),
       .pivot_in   (pivot_in_4_53),
       .start_out  (start_out_4_53),
       .data_out   (data_out_4_53),
       .op_out     (op_out_4_53),
       .pivot_out  (pivot_out_4_53),
       .r          (r_4_53)
     );

  // row 4, col 54

     reg start_in_4_54;
     wire start_out_4_54;

     reg [1:0] op_in_4_54;
     wire [1:0] op_out_4_54;

     wire r_4_54;

     reg data_in_4_54;
     wire data_out_4_54;

     reg pivot_in_4_54;
     wire pivot_out_4_54;

     always @(posedge clk) begin
         op_in_4_54 <= op_out_4_53;
         pivot_in_4_54 <= pivot_out_4_53;
         start_in_4_54 <= start_out_4_53;
     end

     always @(posedge clk) begin
         data_in_4_54 <= data_out_3_54;
     end
  
     processor_AB AB_4_54 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_54),
       .start_in   (start_in_4_54),
       .op_in      (op_in_4_54),
       .pivot_in   (pivot_in_4_54),
       .start_out  (start_out_4_54),
       .data_out   (data_out_4_54),
       .op_out     (op_out_4_54),
       .pivot_out  (pivot_out_4_54),
       .r          (r_4_54)
     );

  // row 4, col 55

     reg start_in_4_55;
     wire start_out_4_55;

     reg [1:0] op_in_4_55;
     wire [1:0] op_out_4_55;

     wire r_4_55;

     reg data_in_4_55;
     wire data_out_4_55;

     reg pivot_in_4_55;
     wire pivot_out_4_55;

     always @(posedge clk) begin
         op_in_4_55 <= op_out_4_54;
         pivot_in_4_55 <= pivot_out_4_54;
         start_in_4_55 <= start_out_4_54;
     end

     always @(posedge clk) begin
         data_in_4_55 <= data_out_3_55;
     end
  
     processor_AB AB_4_55 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_55),
       .start_in   (start_in_4_55),
       .op_in      (op_in_4_55),
       .pivot_in   (pivot_in_4_55),
       .start_out  (start_out_4_55),
       .data_out   (data_out_4_55),
       .op_out     (op_out_4_55),
       .pivot_out  (pivot_out_4_55),
       .r          (r_4_55)
     );

  // row 4, col 56

     reg start_in_4_56;
     wire start_out_4_56;

     reg [1:0] op_in_4_56;
     wire [1:0] op_out_4_56;

     wire r_4_56;

     reg data_in_4_56;
     wire data_out_4_56;

     reg pivot_in_4_56;
     wire pivot_out_4_56;

     always @(posedge clk) begin
         op_in_4_56 <= op_out_4_55;
         pivot_in_4_56 <= pivot_out_4_55;
         start_in_4_56 <= start_out_4_55;
     end

     always @(posedge clk) begin
         data_in_4_56 <= data_out_3_56;
     end
  
     processor_AB AB_4_56 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_56),
       .start_in   (start_in_4_56),
       .op_in      (op_in_4_56),
       .pivot_in   (pivot_in_4_56),
       .start_out  (start_out_4_56),
       .data_out   (data_out_4_56),
       .op_out     (op_out_4_56),
       .pivot_out  (pivot_out_4_56),
       .r          (r_4_56)
     );

  // row 4, col 57

     reg start_in_4_57;
     wire start_out_4_57;

     reg [1:0] op_in_4_57;
     wire [1:0] op_out_4_57;

     wire r_4_57;

     reg data_in_4_57;
     wire data_out_4_57;

     reg pivot_in_4_57;
     wire pivot_out_4_57;

     always @(posedge clk) begin
         op_in_4_57 <= op_out_4_56;
         pivot_in_4_57 <= pivot_out_4_56;
         start_in_4_57 <= start_out_4_56;
     end

     always @(posedge clk) begin
         data_in_4_57 <= data_out_3_57;
     end
  
     processor_AB AB_4_57 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_57),
       .start_in   (start_in_4_57),
       .op_in      (op_in_4_57),
       .pivot_in   (pivot_in_4_57),
       .start_out  (start_out_4_57),
       .data_out   (data_out_4_57),
       .op_out     (op_out_4_57),
       .pivot_out  (pivot_out_4_57),
       .r          (r_4_57)
     );

  // row 4, col 58

     reg start_in_4_58;
     wire start_out_4_58;

     reg [1:0] op_in_4_58;
     wire [1:0] op_out_4_58;

     wire r_4_58;

     reg data_in_4_58;
     wire data_out_4_58;

     reg pivot_in_4_58;
     wire pivot_out_4_58;

     always @(posedge clk) begin
         op_in_4_58 <= op_out_4_57;
         pivot_in_4_58 <= pivot_out_4_57;
         start_in_4_58 <= start_out_4_57;
     end

     always @(posedge clk) begin
         data_in_4_58 <= data_out_3_58;
     end
  
     processor_AB AB_4_58 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_58),
       .start_in   (start_in_4_58),
       .op_in      (op_in_4_58),
       .pivot_in   (pivot_in_4_58),
       .start_out  (start_out_4_58),
       .data_out   (data_out_4_58),
       .op_out     (op_out_4_58),
       .pivot_out  (pivot_out_4_58),
       .r          (r_4_58)
     );

  // row 4, col 59

     reg start_in_4_59;
     wire start_out_4_59;

     reg [1:0] op_in_4_59;
     wire [1:0] op_out_4_59;

     wire r_4_59;

     reg data_in_4_59;
     wire data_out_4_59;

     reg pivot_in_4_59;
     wire pivot_out_4_59;

     always @(posedge clk) begin
         op_in_4_59 <= op_out_4_58;
         pivot_in_4_59 <= pivot_out_4_58;
         start_in_4_59 <= start_out_4_58;
     end

     always @(posedge clk) begin
         data_in_4_59 <= data_out_3_59;
     end
  
     processor_AB AB_4_59 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_59),
       .start_in   (start_in_4_59),
       .op_in      (op_in_4_59),
       .pivot_in   (pivot_in_4_59),
       .start_out  (start_out_4_59),
       .data_out   (data_out_4_59),
       .op_out     (op_out_4_59),
       .pivot_out  (pivot_out_4_59),
       .r          (r_4_59)
     );

  // row 4, col 60

     reg start_in_4_60;
     wire start_out_4_60;

     reg [1:0] op_in_4_60;
     wire [1:0] op_out_4_60;

     wire r_4_60;

     reg data_in_4_60;
     wire data_out_4_60;

     reg pivot_in_4_60;
     wire pivot_out_4_60;

     always @(posedge clk) begin
         op_in_4_60 <= op_out_4_59;
         pivot_in_4_60 <= pivot_out_4_59;
         start_in_4_60 <= start_out_4_59;
     end

     always @(posedge clk) begin
         data_in_4_60 <= data_out_3_60;
     end
  
     processor_AB AB_4_60 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_60),
       .start_in   (start_in_4_60),
       .op_in      (op_in_4_60),
       .pivot_in   (pivot_in_4_60),
       .start_out  (start_out_4_60),
       .data_out   (data_out_4_60),
       .op_out     (op_out_4_60),
       .pivot_out  (pivot_out_4_60),
       .r          (r_4_60)
     );

  // row 4, col 61

     reg start_in_4_61;
     wire start_out_4_61;

     reg [1:0] op_in_4_61;
     wire [1:0] op_out_4_61;

     wire r_4_61;

     reg data_in_4_61;
     wire data_out_4_61;

     reg pivot_in_4_61;
     wire pivot_out_4_61;

     always @(posedge clk) begin
         op_in_4_61 <= op_out_4_60;
         pivot_in_4_61 <= pivot_out_4_60;
         start_in_4_61 <= start_out_4_60;
     end

     always @(posedge clk) begin
         data_in_4_61 <= data_out_3_61;
     end
  
     processor_AB AB_4_61 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_61),
       .start_in   (start_in_4_61),
       .op_in      (op_in_4_61),
       .pivot_in   (pivot_in_4_61),
       .start_out  (start_out_4_61),
       .data_out   (data_out_4_61),
       .op_out     (op_out_4_61),
       .pivot_out  (pivot_out_4_61),
       .r          (r_4_61)
     );

  // row 4, col 62

     reg start_in_4_62;
     wire start_out_4_62;

     reg [1:0] op_in_4_62;
     wire [1:0] op_out_4_62;

     wire r_4_62;

     reg data_in_4_62;
     wire data_out_4_62;

     reg pivot_in_4_62;
     wire pivot_out_4_62;

     always @(posedge clk) begin
         op_in_4_62 <= op_out_4_61;
         pivot_in_4_62 <= pivot_out_4_61;
         start_in_4_62 <= start_out_4_61;
     end

     always @(posedge clk) begin
         data_in_4_62 <= data_out_3_62;
     end
  
     processor_AB AB_4_62 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_62),
       .start_in   (start_in_4_62),
       .op_in      (op_in_4_62),
       .pivot_in   (pivot_in_4_62),
       .start_out  (start_out_4_62),
       .data_out   (data_out_4_62),
       .op_out     (op_out_4_62),
       .pivot_out  (pivot_out_4_62),
       .r          (r_4_62)
     );

  // row 4, col 63

     reg start_in_4_63;
     wire start_out_4_63;

     reg [1:0] op_in_4_63;
     wire [1:0] op_out_4_63;

     wire r_4_63;

     reg data_in_4_63;
     wire data_out_4_63;

     reg pivot_in_4_63;
     wire pivot_out_4_63;

     always @(posedge clk) begin
         op_in_4_63 <= op_out_4_62;
         pivot_in_4_63 <= pivot_out_4_62;
         start_in_4_63 <= start_out_4_62;
     end

     always @(posedge clk) begin
         data_in_4_63 <= data_out_3_63;
     end
  
     processor_AB AB_4_63 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_63),
       .start_in   (start_in_4_63),
       .op_in      (op_in_4_63),
       .pivot_in   (pivot_in_4_63),
       .start_out  (start_out_4_63),
       .data_out   (data_out_4_63),
       .op_out     (op_out_4_63),
       .pivot_out  (pivot_out_4_63),
       .r          (r_4_63)
     );

  // row 4, col 64

     reg start_in_4_64;
     wire start_out_4_64;

     reg [1:0] op_in_4_64;
     wire [1:0] op_out_4_64;

     wire r_4_64;

     reg data_in_4_64;
     wire data_out_4_64;

     reg pivot_in_4_64;
     wire pivot_out_4_64;

     always @(posedge clk) begin
         op_in_4_64 <= op_out_4_63;
         pivot_in_4_64 <= pivot_out_4_63;
         start_in_4_64 <= start_out_4_63;
     end

     always @(posedge clk) begin
         data_in_4_64 <= data_out_3_64;
     end
  
     processor_AB AB_4_64 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_64),
       .start_in   (start_in_4_64),
       .op_in      (op_in_4_64),
       .pivot_in   (pivot_in_4_64),
       .start_out  (start_out_4_64),
       .data_out   (data_out_4_64),
       .op_out     (op_out_4_64),
       .pivot_out  (pivot_out_4_64),
       .r          (r_4_64)
     );

  // row 4, col 65

     reg start_in_4_65;
     wire start_out_4_65;

     reg [1:0] op_in_4_65;
     wire [1:0] op_out_4_65;

     wire r_4_65;

     reg data_in_4_65;
     wire data_out_4_65;

     reg pivot_in_4_65;
     wire pivot_out_4_65;

     always @(posedge clk) begin
         op_in_4_65 <= op_out_4_64;
         pivot_in_4_65 <= pivot_out_4_64;
         start_in_4_65 <= start_out_4_64;
     end

     always @(posedge clk) begin
         data_in_4_65 <= data_out_3_65;
     end
  
     processor_AB AB_4_65 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_65),
       .start_in   (start_in_4_65),
       .op_in      (op_in_4_65),
       .pivot_in   (pivot_in_4_65),
       .start_out  (start_out_4_65),
       .data_out   (data_out_4_65),
       .op_out     (op_out_4_65),
       .pivot_out  (pivot_out_4_65),
       .r          (r_4_65)
     );

  // row 4, col 66

     reg start_in_4_66;
     wire start_out_4_66;

     reg [1:0] op_in_4_66;
     wire [1:0] op_out_4_66;

     wire r_4_66;

     reg data_in_4_66;
     wire data_out_4_66;

     reg pivot_in_4_66;
     wire pivot_out_4_66;

     always @(posedge clk) begin
         op_in_4_66 <= op_out_4_65;
         pivot_in_4_66 <= pivot_out_4_65;
         start_in_4_66 <= start_out_4_65;
     end

     always @(posedge clk) begin
         data_in_4_66 <= data_out_3_66;
     end
  
     processor_AB AB_4_66 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_66),
       .start_in   (start_in_4_66),
       .op_in      (op_in_4_66),
       .pivot_in   (pivot_in_4_66),
       .start_out  (start_out_4_66),
       .data_out   (data_out_4_66),
       .op_out     (op_out_4_66),
       .pivot_out  (pivot_out_4_66),
       .r          (r_4_66)
     );

  // row 4, col 67

     reg start_in_4_67;
     wire start_out_4_67;

     reg [1:0] op_in_4_67;
     wire [1:0] op_out_4_67;

     wire r_4_67;

     reg data_in_4_67;
     wire data_out_4_67;

     reg pivot_in_4_67;
     wire pivot_out_4_67;

     always @(posedge clk) begin
         op_in_4_67 <= op_out_4_66;
         pivot_in_4_67 <= pivot_out_4_66;
         start_in_4_67 <= start_out_4_66;
     end

     always @(posedge clk) begin
         data_in_4_67 <= data_out_3_67;
     end
  
     processor_AB AB_4_67 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_67),
       .start_in   (start_in_4_67),
       .op_in      (op_in_4_67),
       .pivot_in   (pivot_in_4_67),
       .start_out  (start_out_4_67),
       .data_out   (data_out_4_67),
       .op_out     (op_out_4_67),
       .pivot_out  (pivot_out_4_67),
       .r          (r_4_67)
     );

  // row 4, col 68

     reg start_in_4_68;
     wire start_out_4_68;

     reg [1:0] op_in_4_68;
     wire [1:0] op_out_4_68;

     wire r_4_68;

     reg data_in_4_68;
     wire data_out_4_68;

     reg pivot_in_4_68;
     wire pivot_out_4_68;

     always @(posedge clk) begin
         op_in_4_68 <= op_out_4_67;
         pivot_in_4_68 <= pivot_out_4_67;
         start_in_4_68 <= start_out_4_67;
     end

     always @(posedge clk) begin
         data_in_4_68 <= data_out_3_68;
     end
  
     processor_AB AB_4_68 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_68),
       .start_in   (start_in_4_68),
       .op_in      (op_in_4_68),
       .pivot_in   (pivot_in_4_68),
       .start_out  (start_out_4_68),
       .data_out   (data_out_4_68),
       .op_out     (op_out_4_68),
       .pivot_out  (pivot_out_4_68),
       .r          (r_4_68)
     );

  // row 4, col 69

     reg start_in_4_69;
     wire start_out_4_69;

     reg [1:0] op_in_4_69;
     wire [1:0] op_out_4_69;

     wire r_4_69;

     reg data_in_4_69;
     wire data_out_4_69;

     reg pivot_in_4_69;
     wire pivot_out_4_69;

     always @(posedge clk) begin
         op_in_4_69 <= op_out_4_68;
         pivot_in_4_69 <= pivot_out_4_68;
         start_in_4_69 <= start_out_4_68;
     end

     always @(posedge clk) begin
         data_in_4_69 <= data_out_3_69;
     end
  
     processor_AB AB_4_69 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_69),
       .start_in   (start_in_4_69),
       .op_in      (op_in_4_69),
       .pivot_in   (pivot_in_4_69),
       .start_out  (start_out_4_69),
       .data_out   (data_out_4_69),
       .op_out     (op_out_4_69),
       .pivot_out  (pivot_out_4_69),
       .r          (r_4_69)
     );

  // row 4, col 70

     reg start_in_4_70;
     wire start_out_4_70;

     reg [1:0] op_in_4_70;
     wire [1:0] op_out_4_70;

     wire r_4_70;

     reg data_in_4_70;
     wire data_out_4_70;

     reg pivot_in_4_70;
     wire pivot_out_4_70;

     always @(posedge clk) begin
         op_in_4_70 <= op_out_4_69;
         pivot_in_4_70 <= pivot_out_4_69;
         start_in_4_70 <= start_out_4_69;
     end

     always @(posedge clk) begin
         data_in_4_70 <= data_out_3_70;
     end
  
     processor_AB AB_4_70 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_70),
       .start_in   (start_in_4_70),
       .op_in      (op_in_4_70),
       .pivot_in   (pivot_in_4_70),
       .start_out  (start_out_4_70),
       .data_out   (data_out_4_70),
       .op_out     (op_out_4_70),
       .pivot_out  (pivot_out_4_70),
       .r          (r_4_70)
     );

  // row 4, col 71

     reg start_in_4_71;
     wire start_out_4_71;

     reg [1:0] op_in_4_71;
     wire [1:0] op_out_4_71;

     wire r_4_71;

     reg data_in_4_71;
     wire data_out_4_71;

     reg pivot_in_4_71;
     wire pivot_out_4_71;

     always @(posedge clk) begin
         op_in_4_71 <= op_out_4_70;
         pivot_in_4_71 <= pivot_out_4_70;
         start_in_4_71 <= start_out_4_70;
     end

     always @(posedge clk) begin
         data_in_4_71 <= data_out_3_71;
     end
  
     processor_AB AB_4_71 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_71),
       .start_in   (start_in_4_71),
       .op_in      (op_in_4_71),
       .pivot_in   (pivot_in_4_71),
       .start_out  (start_out_4_71),
       .data_out   (data_out_4_71),
       .op_out     (op_out_4_71),
       .pivot_out  (pivot_out_4_71),
       .r          (r_4_71)
     );

  // row 4, col 72

     reg start_in_4_72;
     wire start_out_4_72;

     reg [1:0] op_in_4_72;
     wire [1:0] op_out_4_72;

     wire r_4_72;

     reg data_in_4_72;
     wire data_out_4_72;

     reg pivot_in_4_72;
     wire pivot_out_4_72;

     always @(posedge clk) begin
         op_in_4_72 <= op_out_4_71;
         pivot_in_4_72 <= pivot_out_4_71;
         start_in_4_72 <= start_out_4_71;
     end

     always @(posedge clk) begin
         data_in_4_72 <= data_out_3_72;
     end
  
     processor_AB AB_4_72 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_72),
       .start_in   (start_in_4_72),
       .op_in      (op_in_4_72),
       .pivot_in   (pivot_in_4_72),
       .start_out  (start_out_4_72),
       .data_out   (data_out_4_72),
       .op_out     (op_out_4_72),
       .pivot_out  (pivot_out_4_72),
       .r          (r_4_72)
     );

  // row 4, col 73

     reg start_in_4_73;
     wire start_out_4_73;

     reg [1:0] op_in_4_73;
     wire [1:0] op_out_4_73;

     wire r_4_73;

     reg data_in_4_73;
     wire data_out_4_73;

     reg pivot_in_4_73;
     wire pivot_out_4_73;

     always @(posedge clk) begin
         op_in_4_73 <= op_out_4_72;
         pivot_in_4_73 <= pivot_out_4_72;
         start_in_4_73 <= start_out_4_72;
     end

     always @(posedge clk) begin
         data_in_4_73 <= data_out_3_73;
     end
  
     processor_AB AB_4_73 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_73),
       .start_in   (start_in_4_73),
       .op_in      (op_in_4_73),
       .pivot_in   (pivot_in_4_73),
       .start_out  (start_out_4_73),
       .data_out   (data_out_4_73),
       .op_out     (op_out_4_73),
       .pivot_out  (pivot_out_4_73),
       .r          (r_4_73)
     );

  // row 4, col 74

     reg start_in_4_74;
     wire start_out_4_74;

     reg [1:0] op_in_4_74;
     wire [1:0] op_out_4_74;

     wire r_4_74;

     reg data_in_4_74;
     wire data_out_4_74;

     reg pivot_in_4_74;
     wire pivot_out_4_74;

     always @(posedge clk) begin
         op_in_4_74 <= op_out_4_73;
         pivot_in_4_74 <= pivot_out_4_73;
         start_in_4_74 <= start_out_4_73;
     end

     always @(posedge clk) begin
         data_in_4_74 <= data_out_3_74;
     end
  
     processor_AB AB_4_74 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_74),
       .start_in   (start_in_4_74),
       .op_in      (op_in_4_74),
       .pivot_in   (pivot_in_4_74),
       .start_out  (start_out_4_74),
       .data_out   (data_out_4_74),
       .op_out     (op_out_4_74),
       .pivot_out  (pivot_out_4_74),
       .r          (r_4_74)
     );

  // row 4, col 75

     reg start_in_4_75;
     wire start_out_4_75;

     reg [1:0] op_in_4_75;
     wire [1:0] op_out_4_75;

     wire r_4_75;

     reg data_in_4_75;
     wire data_out_4_75;

     reg pivot_in_4_75;
     wire pivot_out_4_75;

     always @(posedge clk) begin
         op_in_4_75 <= op_out_4_74;
         pivot_in_4_75 <= pivot_out_4_74;
         start_in_4_75 <= start_out_4_74;
     end

     always @(posedge clk) begin
         data_in_4_75 <= data_out_3_75;
     end
  
     processor_AB AB_4_75 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_75),
       .start_in   (start_in_4_75),
       .op_in      (op_in_4_75),
       .pivot_in   (pivot_in_4_75),
       .start_out  (start_out_4_75),
       .data_out   (data_out_4_75),
       .op_out     (op_out_4_75),
       .pivot_out  (pivot_out_4_75),
       .r          (r_4_75)
     );

  // row 4, col 76

     reg start_in_4_76;
     wire start_out_4_76;

     reg [1:0] op_in_4_76;
     wire [1:0] op_out_4_76;

     wire r_4_76;

     reg data_in_4_76;
     wire data_out_4_76;

     reg pivot_in_4_76;
     wire pivot_out_4_76;

     always @(posedge clk) begin
         op_in_4_76 <= op_out_4_75;
         pivot_in_4_76 <= pivot_out_4_75;
         start_in_4_76 <= start_out_4_75;
     end

     always @(posedge clk) begin
         data_in_4_76 <= data_out_3_76;
     end
  
     processor_AB AB_4_76 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_76),
       .start_in   (start_in_4_76),
       .op_in      (op_in_4_76),
       .pivot_in   (pivot_in_4_76),
       .start_out  (start_out_4_76),
       .data_out   (data_out_4_76),
       .op_out     (op_out_4_76),
       .pivot_out  (pivot_out_4_76),
       .r          (r_4_76)
     );

  // row 4, col 77

     reg start_in_4_77;
     wire start_out_4_77;

     reg [1:0] op_in_4_77;
     wire [1:0] op_out_4_77;

     wire r_4_77;

     reg data_in_4_77;
     wire data_out_4_77;

     reg pivot_in_4_77;
     wire pivot_out_4_77;

     always @(posedge clk) begin
         op_in_4_77 <= op_out_4_76;
         pivot_in_4_77 <= pivot_out_4_76;
         start_in_4_77 <= start_out_4_76;
     end

     always @(posedge clk) begin
         data_in_4_77 <= data_out_3_77;
     end
  
     processor_AB AB_4_77 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_77),
       .start_in   (start_in_4_77),
       .op_in      (op_in_4_77),
       .pivot_in   (pivot_in_4_77),
       .start_out  (start_out_4_77),
       .data_out   (data_out_4_77),
       .op_out     (op_out_4_77),
       .pivot_out  (pivot_out_4_77),
       .r          (r_4_77)
     );

  // row 4, col 78

     reg start_in_4_78;
     wire start_out_4_78;

     reg [1:0] op_in_4_78;
     wire [1:0] op_out_4_78;

     wire r_4_78;

     reg data_in_4_78;
     wire data_out_4_78;

     reg pivot_in_4_78;
     wire pivot_out_4_78;

     always @(posedge clk) begin
         op_in_4_78 <= op_out_4_77;
         pivot_in_4_78 <= pivot_out_4_77;
         start_in_4_78 <= start_out_4_77;
     end

     always @(posedge clk) begin
         data_in_4_78 <= data_out_3_78;
     end
  
     processor_AB AB_4_78 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_78),
       .start_in   (start_in_4_78),
       .op_in      (op_in_4_78),
       .pivot_in   (pivot_in_4_78),
       .start_out  (start_out_4_78),
       .data_out   (data_out_4_78),
       .op_out     (op_out_4_78),
       .pivot_out  (pivot_out_4_78),
       .r          (r_4_78)
     );

  // row 4, col 79

     reg start_in_4_79;
     wire start_out_4_79;

     reg [1:0] op_in_4_79;
     wire [1:0] op_out_4_79;

     wire r_4_79;

     reg data_in_4_79;
     wire data_out_4_79;

     reg pivot_in_4_79;
     wire pivot_out_4_79;

     always @(posedge clk) begin
         op_in_4_79 <= op_out_4_78;
         pivot_in_4_79 <= pivot_out_4_78;
         start_in_4_79 <= start_out_4_78;
     end

     always @(posedge clk) begin
         data_in_4_79 <= data_out_3_79;
     end
  
     processor_AB AB_4_79 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_79),
       .start_in   (start_in_4_79),
       .op_in      (op_in_4_79),
       .pivot_in   (pivot_in_4_79),
       .start_out  (start_out_4_79),
       .data_out   (data_out_4_79),
       .op_out     (op_out_4_79),
       .pivot_out  (pivot_out_4_79),
       .r          (r_4_79)
     );

  // row 4, col 80

     reg start_in_4_80;
     wire start_out_4_80;

     reg [1:0] op_in_4_80;
     wire [1:0] op_out_4_80;

     wire r_4_80;

     reg data_in_4_80;
     wire data_out_4_80;

     reg pivot_in_4_80;
     wire pivot_out_4_80;

     always @(posedge clk) begin
         op_in_4_80 <= op_out_4_79;
         pivot_in_4_80 <= pivot_out_4_79;
         start_in_4_80 <= start_out_4_79;
     end

     always @(posedge clk) begin
         data_in_4_80 <= data_out_3_80;
     end
  
     processor_AB AB_4_80 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_80),
       .start_in   (start_in_4_80),
       .op_in      (op_in_4_80),
       .pivot_in   (pivot_in_4_80),
       .start_out  (start_out_4_80),
       .data_out   (data_out_4_80),
       .op_out     (op_out_4_80),
       .pivot_out  (pivot_out_4_80),
       .r          (r_4_80)
     );

  // row 4, col 81

     reg start_in_4_81;
     wire start_out_4_81;

     reg [1:0] op_in_4_81;
     wire [1:0] op_out_4_81;

     wire r_4_81;

     reg data_in_4_81;
     wire data_out_4_81;

     reg pivot_in_4_81;
     wire pivot_out_4_81;

     always @(posedge clk) begin
         op_in_4_81 <= op_out_4_80;
         pivot_in_4_81 <= pivot_out_4_80;
         start_in_4_81 <= start_out_4_80;
     end

     always @(posedge clk) begin
         data_in_4_81 <= data_out_3_81;
     end
  
     processor_AB AB_4_81 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_81),
       .start_in   (start_in_4_81),
       .op_in      (op_in_4_81),
       .pivot_in   (pivot_in_4_81),
       .start_out  (start_out_4_81),
       .data_out   (data_out_4_81),
       .op_out     (op_out_4_81),
       .pivot_out  (pivot_out_4_81),
       .r          (r_4_81)
     );

  // row 4, col 82

     reg start_in_4_82;
     wire start_out_4_82;

     reg [1:0] op_in_4_82;
     wire [1:0] op_out_4_82;

     wire r_4_82;

     reg data_in_4_82;
     wire data_out_4_82;

     reg pivot_in_4_82;
     wire pivot_out_4_82;

     always @(posedge clk) begin
         op_in_4_82 <= op_out_4_81;
         pivot_in_4_82 <= pivot_out_4_81;
         start_in_4_82 <= start_out_4_81;
     end

     always @(posedge clk) begin
         data_in_4_82 <= data_out_3_82;
     end
  
     processor_AB AB_4_82 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_82),
       .start_in   (start_in_4_82),
       .op_in      (op_in_4_82),
       .pivot_in   (pivot_in_4_82),
       .start_out  (start_out_4_82),
       .data_out   (data_out_4_82),
       .op_out     (op_out_4_82),
       .pivot_out  (pivot_out_4_82),
       .r          (r_4_82)
     );

  // row 4, col 83

     reg start_in_4_83;
     wire start_out_4_83;

     reg [1:0] op_in_4_83;
     wire [1:0] op_out_4_83;

     wire r_4_83;

     reg data_in_4_83;
     wire data_out_4_83;

     reg pivot_in_4_83;
     wire pivot_out_4_83;

     always @(posedge clk) begin
         op_in_4_83 <= op_out_4_82;
         pivot_in_4_83 <= pivot_out_4_82;
         start_in_4_83 <= start_out_4_82;
     end

     always @(posedge clk) begin
         data_in_4_83 <= data_out_3_83;
     end
  
     processor_AB AB_4_83 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_83),
       .start_in   (start_in_4_83),
       .op_in      (op_in_4_83),
       .pivot_in   (pivot_in_4_83),
       .start_out  (start_out_4_83),
       .data_out   (data_out_4_83),
       .op_out     (op_out_4_83),
       .pivot_out  (pivot_out_4_83),
       .r          (r_4_83)
     );

  // row 4, col 84

     reg start_in_4_84;
     wire start_out_4_84;

     reg [1:0] op_in_4_84;
     wire [1:0] op_out_4_84;

     wire r_4_84;

     reg data_in_4_84;
     wire data_out_4_84;

     reg pivot_in_4_84;
     wire pivot_out_4_84;

     always @(posedge clk) begin
         op_in_4_84 <= op_out_4_83;
         pivot_in_4_84 <= pivot_out_4_83;
         start_in_4_84 <= start_out_4_83;
     end

     always @(posedge clk) begin
         data_in_4_84 <= data_out_3_84;
     end
  
     processor_AB AB_4_84 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_84),
       .start_in   (start_in_4_84),
       .op_in      (op_in_4_84),
       .pivot_in   (pivot_in_4_84),
       .start_out  (start_out_4_84),
       .data_out   (data_out_4_84),
       .op_out     (op_out_4_84),
       .pivot_out  (pivot_out_4_84),
       .r          (r_4_84)
     );

  // row 4, col 85

     reg start_in_4_85;
     wire start_out_4_85;

     reg [1:0] op_in_4_85;
     wire [1:0] op_out_4_85;

     wire r_4_85;

     reg data_in_4_85;
     wire data_out_4_85;

     reg pivot_in_4_85;
     wire pivot_out_4_85;

     always @(posedge clk) begin
         op_in_4_85 <= op_out_4_84;
         pivot_in_4_85 <= pivot_out_4_84;
         start_in_4_85 <= start_out_4_84;
     end

     always @(posedge clk) begin
         data_in_4_85 <= data_out_3_85;
     end
  
     processor_AB AB_4_85 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_85),
       .start_in   (start_in_4_85),
       .op_in      (op_in_4_85),
       .pivot_in   (pivot_in_4_85),
       .start_out  (start_out_4_85),
       .data_out   (data_out_4_85),
       .op_out     (op_out_4_85),
       .pivot_out  (pivot_out_4_85),
       .r          (r_4_85)
     );

  // row 4, col 86

     reg start_in_4_86;
     wire start_out_4_86;

     reg [1:0] op_in_4_86;
     wire [1:0] op_out_4_86;

     wire r_4_86;

     reg data_in_4_86;
     wire data_out_4_86;

     reg pivot_in_4_86;
     wire pivot_out_4_86;

     always @(posedge clk) begin
         op_in_4_86 <= op_out_4_85;
         pivot_in_4_86 <= pivot_out_4_85;
         start_in_4_86 <= start_out_4_85;
     end

     always @(posedge clk) begin
         data_in_4_86 <= data_out_3_86;
     end
  
     processor_AB AB_4_86 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_86),
       .start_in   (start_in_4_86),
       .op_in      (op_in_4_86),
       .pivot_in   (pivot_in_4_86),
       .start_out  (start_out_4_86),
       .data_out   (data_out_4_86),
       .op_out     (op_out_4_86),
       .pivot_out  (pivot_out_4_86),
       .r          (r_4_86)
     );

  // row 4, col 87

     reg start_in_4_87;
     wire start_out_4_87;

     reg [1:0] op_in_4_87;
     wire [1:0] op_out_4_87;

     wire r_4_87;

     reg data_in_4_87;
     wire data_out_4_87;

     reg pivot_in_4_87;
     wire pivot_out_4_87;

     always @(posedge clk) begin
         op_in_4_87 <= op_out_4_86;
         pivot_in_4_87 <= pivot_out_4_86;
         start_in_4_87 <= start_out_4_86;
     end

     always @(posedge clk) begin
         data_in_4_87 <= data_out_3_87;
     end
  
     processor_AB AB_4_87 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_87),
       .start_in   (start_in_4_87),
       .op_in      (op_in_4_87),
       .pivot_in   (pivot_in_4_87),
       .start_out  (start_out_4_87),
       .data_out   (data_out_4_87),
       .op_out     (op_out_4_87),
       .pivot_out  (pivot_out_4_87),
       .r          (r_4_87)
     );

  // row 4, col 88

     reg start_in_4_88;
     wire start_out_4_88;

     reg [1:0] op_in_4_88;
     wire [1:0] op_out_4_88;

     wire r_4_88;

     reg data_in_4_88;
     wire data_out_4_88;

     reg pivot_in_4_88;
     wire pivot_out_4_88;

     always @(posedge clk) begin
         op_in_4_88 <= op_out_4_87;
         pivot_in_4_88 <= pivot_out_4_87;
         start_in_4_88 <= start_out_4_87;
     end

     always @(posedge clk) begin
         data_in_4_88 <= data_out_3_88;
     end
  
     processor_AB AB_4_88 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_88),
       .start_in   (start_in_4_88),
       .op_in      (op_in_4_88),
       .pivot_in   (pivot_in_4_88),
       .start_out  (start_out_4_88),
       .data_out   (data_out_4_88),
       .op_out     (op_out_4_88),
       .pivot_out  (pivot_out_4_88),
       .r          (r_4_88)
     );

  // row 4, col 89

     reg start_in_4_89;
     wire start_out_4_89;

     reg [1:0] op_in_4_89;
     wire [1:0] op_out_4_89;

     wire r_4_89;

     reg data_in_4_89;
     wire data_out_4_89;

     reg pivot_in_4_89;
     wire pivot_out_4_89;

     always @(posedge clk) begin
         op_in_4_89 <= op_out_4_88;
         pivot_in_4_89 <= pivot_out_4_88;
         start_in_4_89 <= start_out_4_88;
     end

     always @(posedge clk) begin
         data_in_4_89 <= data_out_3_89;
     end
  
     processor_AB AB_4_89 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_89),
       .start_in   (start_in_4_89),
       .op_in      (op_in_4_89),
       .pivot_in   (pivot_in_4_89),
       .start_out  (start_out_4_89),
       .data_out   (data_out_4_89),
       .op_out     (op_out_4_89),
       .pivot_out  (pivot_out_4_89),
       .r          (r_4_89)
     );

  // row 4, col 90

     reg start_in_4_90;
     wire start_out_4_90;

     reg [1:0] op_in_4_90;
     wire [1:0] op_out_4_90;

     wire r_4_90;

     reg data_in_4_90;
     wire data_out_4_90;

     reg pivot_in_4_90;
     wire pivot_out_4_90;

     always @(posedge clk) begin
         op_in_4_90 <= op_out_4_89;
         pivot_in_4_90 <= pivot_out_4_89;
         start_in_4_90 <= start_out_4_89;
     end

     always @(posedge clk) begin
         data_in_4_90 <= data_out_3_90;
     end
  
     processor_AB AB_4_90 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_90),
       .start_in   (start_in_4_90),
       .op_in      (op_in_4_90),
       .pivot_in   (pivot_in_4_90),
       .start_out  (start_out_4_90),
       .data_out   (data_out_4_90),
       .op_out     (op_out_4_90),
       .pivot_out  (pivot_out_4_90),
       .r          (r_4_90)
     );

  // row 4, col 91

     reg start_in_4_91;
     wire start_out_4_91;

     reg [1:0] op_in_4_91;
     wire [1:0] op_out_4_91;

     wire r_4_91;

     reg data_in_4_91;
     wire data_out_4_91;

     reg pivot_in_4_91;
     wire pivot_out_4_91;

     always @(posedge clk) begin
         op_in_4_91 <= op_out_4_90;
         pivot_in_4_91 <= pivot_out_4_90;
         start_in_4_91 <= start_out_4_90;
     end

     always @(posedge clk) begin
         data_in_4_91 <= data_out_3_91;
     end
  
     processor_AB AB_4_91 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_91),
       .start_in   (start_in_4_91),
       .op_in      (op_in_4_91),
       .pivot_in   (pivot_in_4_91),
       .start_out  (start_out_4_91),
       .data_out   (data_out_4_91),
       .op_out     (op_out_4_91),
       .pivot_out  (pivot_out_4_91),
       .r          (r_4_91)
     );

  // row 4, col 92

     reg start_in_4_92;
     wire start_out_4_92;

     reg [1:0] op_in_4_92;
     wire [1:0] op_out_4_92;

     wire r_4_92;

     reg data_in_4_92;
     wire data_out_4_92;

     reg pivot_in_4_92;
     wire pivot_out_4_92;

     always @(posedge clk) begin
         op_in_4_92 <= op_out_4_91;
         pivot_in_4_92 <= pivot_out_4_91;
         start_in_4_92 <= start_out_4_91;
     end

     always @(posedge clk) begin
         data_in_4_92 <= data_out_3_92;
     end
  
     processor_AB AB_4_92 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_92),
       .start_in   (start_in_4_92),
       .op_in      (op_in_4_92),
       .pivot_in   (pivot_in_4_92),
       .start_out  (start_out_4_92),
       .data_out   (data_out_4_92),
       .op_out     (op_out_4_92),
       .pivot_out  (pivot_out_4_92),
       .r          (r_4_92)
     );

  // row 4, col 93

     reg start_in_4_93;
     wire start_out_4_93;

     reg [1:0] op_in_4_93;
     wire [1:0] op_out_4_93;

     wire r_4_93;

     reg data_in_4_93;
     wire data_out_4_93;

     reg pivot_in_4_93;
     wire pivot_out_4_93;

     always @(posedge clk) begin
         op_in_4_93 <= op_out_4_92;
         pivot_in_4_93 <= pivot_out_4_92;
         start_in_4_93 <= start_out_4_92;
     end

     always @(posedge clk) begin
         data_in_4_93 <= data_out_3_93;
     end
  
     processor_AB AB_4_93 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_93),
       .start_in   (start_in_4_93),
       .op_in      (op_in_4_93),
       .pivot_in   (pivot_in_4_93),
       .start_out  (start_out_4_93),
       .data_out   (data_out_4_93),
       .op_out     (op_out_4_93),
       .pivot_out  (pivot_out_4_93),
       .r          (r_4_93)
     );

  // row 4, col 94

     reg start_in_4_94;
     wire start_out_4_94;

     reg [1:0] op_in_4_94;
     wire [1:0] op_out_4_94;

     wire r_4_94;

     reg data_in_4_94;
     wire data_out_4_94;

     reg pivot_in_4_94;
     wire pivot_out_4_94;

     always @(posedge clk) begin
         op_in_4_94 <= op_out_4_93;
         pivot_in_4_94 <= pivot_out_4_93;
         start_in_4_94 <= start_out_4_93;
     end

     always @(posedge clk) begin
         data_in_4_94 <= data_out_3_94;
     end
  
     processor_AB AB_4_94 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_94),
       .start_in   (start_in_4_94),
       .op_in      (op_in_4_94),
       .pivot_in   (pivot_in_4_94),
       .start_out  (start_out_4_94),
       .data_out   (data_out_4_94),
       .op_out     (op_out_4_94),
       .pivot_out  (pivot_out_4_94),
       .r          (r_4_94)
     );

  // row 4, col 95

     reg start_in_4_95;
     wire start_out_4_95;

     reg [1:0] op_in_4_95;
     wire [1:0] op_out_4_95;

     wire r_4_95;

     reg data_in_4_95;
     wire data_out_4_95;

     reg pivot_in_4_95;
     wire pivot_out_4_95;

     always @(posedge clk) begin
         op_in_4_95 <= op_out_4_94;
         pivot_in_4_95 <= pivot_out_4_94;
         start_in_4_95 <= start_out_4_94;
     end

     always @(posedge clk) begin
         data_in_4_95 <= data_out_3_95;
     end
  
     processor_AB AB_4_95 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_95),
       .start_in   (start_in_4_95),
       .op_in      (op_in_4_95),
       .pivot_in   (pivot_in_4_95),
       .start_out  (start_out_4_95),
       .data_out   (data_out_4_95),
       .op_out     (op_out_4_95),
       .pivot_out  (pivot_out_4_95),
       .r          (r_4_95)
     );

  // row 4, col 96

     reg start_in_4_96;
     wire start_out_4_96;

     reg [1:0] op_in_4_96;
     wire [1:0] op_out_4_96;

     wire r_4_96;

     reg data_in_4_96;
     wire data_out_4_96;

     reg pivot_in_4_96;
     wire pivot_out_4_96;

     always @(posedge clk) begin
         op_in_4_96 <= op_out_4_95;
         pivot_in_4_96 <= pivot_out_4_95;
         start_in_4_96 <= start_out_4_95;
     end

     always @(posedge clk) begin
         data_in_4_96 <= data_out_3_96;
     end
  
     processor_AB AB_4_96 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_96),
       .start_in   (start_in_4_96),
       .op_in      (op_in_4_96),
       .pivot_in   (pivot_in_4_96),
       .start_out  (start_out_4_96),
       .data_out   (data_out_4_96),
       .op_out     (op_out_4_96),
       .pivot_out  (pivot_out_4_96),
       .r          (r_4_96)
     );

  // row 4, col 97

     reg start_in_4_97;
     wire start_out_4_97;

     reg [1:0] op_in_4_97;
     wire [1:0] op_out_4_97;

     wire r_4_97;

     reg data_in_4_97;
     wire data_out_4_97;

     reg pivot_in_4_97;
     wire pivot_out_4_97;

     always @(posedge clk) begin
         op_in_4_97 <= op_out_4_96;
         pivot_in_4_97 <= pivot_out_4_96;
         start_in_4_97 <= start_out_4_96;
     end

     always @(posedge clk) begin
         data_in_4_97 <= data_out_3_97;
     end
  
     processor_AB AB_4_97 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_97),
       .start_in   (start_in_4_97),
       .op_in      (op_in_4_97),
       .pivot_in   (pivot_in_4_97),
       .start_out  (start_out_4_97),
       .data_out   (data_out_4_97),
       .op_out     (op_out_4_97),
       .pivot_out  (pivot_out_4_97),
       .r          (r_4_97)
     );

  // row 4, col 98

     reg start_in_4_98;
     wire start_out_4_98;

     reg [1:0] op_in_4_98;
     wire [1:0] op_out_4_98;

     wire r_4_98;

     reg data_in_4_98;
     wire data_out_4_98;

     reg pivot_in_4_98;
     wire pivot_out_4_98;

     always @(posedge clk) begin
         op_in_4_98 <= op_out_4_97;
         pivot_in_4_98 <= pivot_out_4_97;
         start_in_4_98 <= start_out_4_97;
     end

     always @(posedge clk) begin
         data_in_4_98 <= data_out_3_98;
     end
  
     processor_AB AB_4_98 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_98),
       .start_in   (start_in_4_98),
       .op_in      (op_in_4_98),
       .pivot_in   (pivot_in_4_98),
       .start_out  (start_out_4_98),
       .data_out   (data_out_4_98),
       .op_out     (op_out_4_98),
       .pivot_out  (pivot_out_4_98),
       .r          (r_4_98)
     );

  // row 4, col 99

     reg start_in_4_99;
     wire start_out_4_99;

     reg [1:0] op_in_4_99;
     wire [1:0] op_out_4_99;

     wire r_4_99;

     reg data_in_4_99;
     wire data_out_4_99;

     reg pivot_in_4_99;
     wire pivot_out_4_99;

     always @(posedge clk) begin
         op_in_4_99 <= op_out_4_98;
         pivot_in_4_99 <= pivot_out_4_98;
         start_in_4_99 <= start_out_4_98;
     end

     always @(posedge clk) begin
         data_in_4_99 <= data_out_3_99;
     end
  
     processor_AB AB_4_99 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_99),
       .start_in   (start_in_4_99),
       .op_in      (op_in_4_99),
       .pivot_in   (pivot_in_4_99),
       .start_out  (start_out_4_99),
       .data_out   (data_out_4_99),
       .op_out     (op_out_4_99),
       .pivot_out  (pivot_out_4_99),
       .r          (r_4_99)
     );

  // row 4, col 100

     reg start_in_4_100;
     wire start_out_4_100;

     reg [1:0] op_in_4_100;
     wire [1:0] op_out_4_100;

     wire r_4_100;

     reg data_in_4_100;
     wire data_out_4_100;

     reg pivot_in_4_100;
     wire pivot_out_4_100;

     always @(posedge clk) begin
         op_in_4_100 <= op_out_4_99;
         pivot_in_4_100 <= pivot_out_4_99;
         start_in_4_100 <= start_out_4_99;
     end

     always @(posedge clk) begin
         data_in_4_100 <= data_out_3_100;
     end
  
     processor_AB AB_4_100 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_100),
       .start_in   (start_in_4_100),
       .op_in      (op_in_4_100),
       .pivot_in   (pivot_in_4_100),
       .start_out  (start_out_4_100),
       .data_out   (data_out_4_100),
       .op_out     (op_out_4_100),
       .pivot_out  (pivot_out_4_100),
       .r          (r_4_100)
     );

  /////////////////////////////////////
  // row 5
  // row 5, col 0

     wire start_in_5_0;
     wire start_out_5_0;

     wire [1:0] op_in_5_0;
     wire [1:0] op_out_5_0;

     wire r_5_0;

     reg data_in_5_0;
     wire data_out_5_0;

     wire pivot_in_5_0;
     wire pivout_out_5_0;

     assign op_in_5_0 = mode & start ? 2'b01 : 2'b00;
     assign pivot_in_5_0 = 0;

     assign start_in_5_0 = start_row[5]; 

     always @(posedge clk) begin
         data_in_5_0 <= data_out_4_0;
     end

     processor_AB AB_5_0 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_0),
       .start_in   (start_in_5_0),
       .op_in      (op_in_5_0),
       .pivot_in   (pivot_in_5_0),
       .start_out  (start_out_5_0),
       .data_out   (data_out_5_0),
       .op_out     (op_out_5_0),
       .pivot_out  (pivot_out_5_0),
       .r          (r_5_0)
     );

  // row 5, col 1

     reg start_in_5_1;
     wire start_out_5_1;

     reg [1:0] op_in_5_1;
     wire [1:0] op_out_5_1;

     wire r_5_1;

     reg data_in_5_1;
     wire data_out_5_1;

     reg pivot_in_5_1;
     wire pivot_out_5_1;

     always @(posedge clk) begin
         op_in_5_1 <= op_out_5_0;
         pivot_in_5_1 <= pivot_out_5_0;
         start_in_5_1 <= start_out_5_0;
     end

     always @(posedge clk) begin
         data_in_5_1 <= data_out_4_1;
     end
  
     processor_AB AB_5_1 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_1),
       .start_in   (start_in_5_1),
       .op_in      (op_in_5_1),
       .pivot_in   (pivot_in_5_1),
       .start_out  (start_out_5_1),
       .data_out   (data_out_5_1),
       .op_out     (op_out_5_1),
       .pivot_out  (pivot_out_5_1),
       .r          (r_5_1)
     );

  // row 5, col 2

     reg start_in_5_2;
     wire start_out_5_2;

     reg [1:0] op_in_5_2;
     wire [1:0] op_out_5_2;

     wire r_5_2;

     reg data_in_5_2;
     wire data_out_5_2;

     reg pivot_in_5_2;
     wire pivot_out_5_2;

     always @(posedge clk) begin
         op_in_5_2 <= op_out_5_1;
         pivot_in_5_2 <= pivot_out_5_1;
         start_in_5_2 <= start_out_5_1;
     end

     always @(posedge clk) begin
         data_in_5_2 <= data_out_4_2;
     end
  
     processor_AB AB_5_2 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_2),
       .start_in   (start_in_5_2),
       .op_in      (op_in_5_2),
       .pivot_in   (pivot_in_5_2),
       .start_out  (start_out_5_2),
       .data_out   (data_out_5_2),
       .op_out     (op_out_5_2),
       .pivot_out  (pivot_out_5_2),
       .r          (r_5_2)
     );

  // row 5, col 3

     reg start_in_5_3;
     wire start_out_5_3;

     reg [1:0] op_in_5_3;
     wire [1:0] op_out_5_3;

     wire r_5_3;

     reg data_in_5_3;
     wire data_out_5_3;

     reg pivot_in_5_3;
     wire pivot_out_5_3;

     always @(posedge clk) begin
         op_in_5_3 <= op_out_5_2;
         pivot_in_5_3 <= pivot_out_5_2;
         start_in_5_3 <= start_out_5_2;
     end

     always @(posedge clk) begin
         data_in_5_3 <= data_out_4_3;
     end
  
     processor_AB AB_5_3 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_3),
       .start_in   (start_in_5_3),
       .op_in      (op_in_5_3),
       .pivot_in   (pivot_in_5_3),
       .start_out  (start_out_5_3),
       .data_out   (data_out_5_3),
       .op_out     (op_out_5_3),
       .pivot_out  (pivot_out_5_3),
       .r          (r_5_3)
     );

  // row 5, col 4

     reg start_in_5_4;
     wire start_out_5_4;

     reg [1:0] op_in_5_4;
     wire [1:0] op_out_5_4;

     wire r_5_4;

     reg data_in_5_4;
     wire data_out_5_4;

     reg pivot_in_5_4;
     wire pivot_out_5_4;

     always @(posedge clk) begin
         op_in_5_4 <= op_out_5_3;
         pivot_in_5_4 <= pivot_out_5_3;
         start_in_5_4 <= start_out_5_3;
     end

     always @(posedge clk) begin
         data_in_5_4 <= data_out_4_4;
     end
  
     processor_AB AB_5_4 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_4),
       .start_in   (start_in_5_4),
       .op_in      (op_in_5_4),
       .pivot_in   (pivot_in_5_4),
       .start_out  (start_out_5_4),
       .data_out   (data_out_5_4),
       .op_out     (op_out_5_4),
       .pivot_out  (pivot_out_5_4),
       .r          (r_5_4)
     );

  // row 5, col 5

     reg start_in_5_5;
     wire start_out_5_5;

     reg [1:0] op_in_5_5;
     wire [1:0] op_out_5_5;

     wire r_5_5;

     reg data_in_5_5;
     wire data_out_5_5;

     reg pivot_in_5_5;
     wire pivot_out_5_5;

     always @(posedge clk) begin
         op_in_5_5 <= op_out_5_4;
         pivot_in_5_5 <= pivot_out_5_4;
         start_in_5_5 <= start_out_5_4;
     end

     always @(posedge clk) begin
         data_in_5_5 <= data_out_4_5;
     end
  
     processor_AB AB_5_5 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_5),
       .start_in   (start_in_5_5),
       .op_in      (op_in_5_5),
       .pivot_in   (pivot_in_5_5),
       .start_out  (start_out_5_5),
       .data_out   (data_out_5_5),
       .op_out     (op_out_5_5),
       .pivot_out  (pivot_out_5_5),
       .r          (r_5_5)
     );

  // row 5, col 6

     reg start_in_5_6;
     wire start_out_5_6;

     reg [1:0] op_in_5_6;
     wire [1:0] op_out_5_6;

     wire r_5_6;

     reg data_in_5_6;
     wire data_out_5_6;

     reg pivot_in_5_6;
     wire pivot_out_5_6;

     always @(posedge clk) begin
         op_in_5_6 <= op_out_5_5;
         pivot_in_5_6 <= pivot_out_5_5;
         start_in_5_6 <= start_out_5_5;
     end

     always @(posedge clk) begin
         data_in_5_6 <= data_out_4_6;
     end
  
     processor_AB AB_5_6 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_6),
       .start_in   (start_in_5_6),
       .op_in      (op_in_5_6),
       .pivot_in   (pivot_in_5_6),
       .start_out  (start_out_5_6),
       .data_out   (data_out_5_6),
       .op_out     (op_out_5_6),
       .pivot_out  (pivot_out_5_6),
       .r          (r_5_6)
     );

  // row 5, col 7

     reg start_in_5_7;
     wire start_out_5_7;

     reg [1:0] op_in_5_7;
     wire [1:0] op_out_5_7;

     wire r_5_7;

     reg data_in_5_7;
     wire data_out_5_7;

     reg pivot_in_5_7;
     wire pivot_out_5_7;

     always @(posedge clk) begin
         op_in_5_7 <= op_out_5_6;
         pivot_in_5_7 <= pivot_out_5_6;
         start_in_5_7 <= start_out_5_6;
     end

     always @(posedge clk) begin
         data_in_5_7 <= data_out_4_7;
     end
  
     processor_AB AB_5_7 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_7),
       .start_in   (start_in_5_7),
       .op_in      (op_in_5_7),
       .pivot_in   (pivot_in_5_7),
       .start_out  (start_out_5_7),
       .data_out   (data_out_5_7),
       .op_out     (op_out_5_7),
       .pivot_out  (pivot_out_5_7),
       .r          (r_5_7)
     );

  // row 5, col 8

     reg start_in_5_8;
     wire start_out_5_8;

     reg [1:0] op_in_5_8;
     wire [1:0] op_out_5_8;

     wire r_5_8;

     reg data_in_5_8;
     wire data_out_5_8;

     reg pivot_in_5_8;
     wire pivot_out_5_8;

     always @(posedge clk) begin
         op_in_5_8 <= op_out_5_7;
         pivot_in_5_8 <= pivot_out_5_7;
         start_in_5_8 <= start_out_5_7;
     end

     always @(posedge clk) begin
         data_in_5_8 <= data_out_4_8;
     end
  
     processor_AB AB_5_8 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_8),
       .start_in   (start_in_5_8),
       .op_in      (op_in_5_8),
       .pivot_in   (pivot_in_5_8),
       .start_out  (start_out_5_8),
       .data_out   (data_out_5_8),
       .op_out     (op_out_5_8),
       .pivot_out  (pivot_out_5_8),
       .r          (r_5_8)
     );

  // row 5, col 9

     reg start_in_5_9;
     wire start_out_5_9;

     reg [1:0] op_in_5_9;
     wire [1:0] op_out_5_9;

     wire r_5_9;

     reg data_in_5_9;
     wire data_out_5_9;

     reg pivot_in_5_9;
     wire pivot_out_5_9;

     always @(posedge clk) begin
         op_in_5_9 <= op_out_5_8;
         pivot_in_5_9 <= pivot_out_5_8;
         start_in_5_9 <= start_out_5_8;
     end

     always @(posedge clk) begin
         data_in_5_9 <= data_out_4_9;
     end
  
     processor_AB AB_5_9 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_9),
       .start_in   (start_in_5_9),
       .op_in      (op_in_5_9),
       .pivot_in   (pivot_in_5_9),
       .start_out  (start_out_5_9),
       .data_out   (data_out_5_9),
       .op_out     (op_out_5_9),
       .pivot_out  (pivot_out_5_9),
       .r          (r_5_9)
     );

  // row 5, col 10

     reg start_in_5_10;
     wire start_out_5_10;

     reg [1:0] op_in_5_10;
     wire [1:0] op_out_5_10;

     wire r_5_10;

     reg data_in_5_10;
     wire data_out_5_10;

     reg pivot_in_5_10;
     wire pivot_out_5_10;

     always @(posedge clk) begin
         op_in_5_10 <= op_out_5_9;
         pivot_in_5_10 <= pivot_out_5_9;
         start_in_5_10 <= start_out_5_9;
     end

     always @(posedge clk) begin
         data_in_5_10 <= data_out_4_10;
     end
  
     processor_AB AB_5_10 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_10),
       .start_in   (start_in_5_10),
       .op_in      (op_in_5_10),
       .pivot_in   (pivot_in_5_10),
       .start_out  (start_out_5_10),
       .data_out   (data_out_5_10),
       .op_out     (op_out_5_10),
       .pivot_out  (pivot_out_5_10),
       .r          (r_5_10)
     );

  // row 5, col 11

     reg start_in_5_11;
     wire start_out_5_11;

     reg [1:0] op_in_5_11;
     wire [1:0] op_out_5_11;

     wire r_5_11;

     reg data_in_5_11;
     wire data_out_5_11;

     reg pivot_in_5_11;
     wire pivot_out_5_11;

     always @(posedge clk) begin
         op_in_5_11 <= op_out_5_10;
         pivot_in_5_11 <= pivot_out_5_10;
         start_in_5_11 <= start_out_5_10;
     end

     always @(posedge clk) begin
         data_in_5_11 <= data_out_4_11;
     end
  
     processor_AB AB_5_11 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_11),
       .start_in   (start_in_5_11),
       .op_in      (op_in_5_11),
       .pivot_in   (pivot_in_5_11),
       .start_out  (start_out_5_11),
       .data_out   (data_out_5_11),
       .op_out     (op_out_5_11),
       .pivot_out  (pivot_out_5_11),
       .r          (r_5_11)
     );

  // row 5, col 12

     reg start_in_5_12;
     wire start_out_5_12;

     reg [1:0] op_in_5_12;
     wire [1:0] op_out_5_12;

     wire r_5_12;

     reg data_in_5_12;
     wire data_out_5_12;

     reg pivot_in_5_12;
     wire pivot_out_5_12;

     always @(posedge clk) begin
         op_in_5_12 <= op_out_5_11;
         pivot_in_5_12 <= pivot_out_5_11;
         start_in_5_12 <= start_out_5_11;
     end

     always @(posedge clk) begin
         data_in_5_12 <= data_out_4_12;
     end
  
     processor_AB AB_5_12 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_12),
       .start_in   (start_in_5_12),
       .op_in      (op_in_5_12),
       .pivot_in   (pivot_in_5_12),
       .start_out  (start_out_5_12),
       .data_out   (data_out_5_12),
       .op_out     (op_out_5_12),
       .pivot_out  (pivot_out_5_12),
       .r          (r_5_12)
     );

  // row 5, col 13

     reg start_in_5_13;
     wire start_out_5_13;

     reg [1:0] op_in_5_13;
     wire [1:0] op_out_5_13;

     wire r_5_13;

     reg data_in_5_13;
     wire data_out_5_13;

     reg pivot_in_5_13;
     wire pivot_out_5_13;

     always @(posedge clk) begin
         op_in_5_13 <= op_out_5_12;
         pivot_in_5_13 <= pivot_out_5_12;
         start_in_5_13 <= start_out_5_12;
     end

     always @(posedge clk) begin
         data_in_5_13 <= data_out_4_13;
     end
  
     processor_AB AB_5_13 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_13),
       .start_in   (start_in_5_13),
       .op_in      (op_in_5_13),
       .pivot_in   (pivot_in_5_13),
       .start_out  (start_out_5_13),
       .data_out   (data_out_5_13),
       .op_out     (op_out_5_13),
       .pivot_out  (pivot_out_5_13),
       .r          (r_5_13)
     );

  // row 5, col 14

     reg start_in_5_14;
     wire start_out_5_14;

     reg [1:0] op_in_5_14;
     wire [1:0] op_out_5_14;

     wire r_5_14;

     reg data_in_5_14;
     wire data_out_5_14;

     reg pivot_in_5_14;
     wire pivot_out_5_14;

     always @(posedge clk) begin
         op_in_5_14 <= op_out_5_13;
         pivot_in_5_14 <= pivot_out_5_13;
         start_in_5_14 <= start_out_5_13;
     end

     always @(posedge clk) begin
         data_in_5_14 <= data_out_4_14;
     end
  
     processor_AB AB_5_14 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_14),
       .start_in   (start_in_5_14),
       .op_in      (op_in_5_14),
       .pivot_in   (pivot_in_5_14),
       .start_out  (start_out_5_14),
       .data_out   (data_out_5_14),
       .op_out     (op_out_5_14),
       .pivot_out  (pivot_out_5_14),
       .r          (r_5_14)
     );

  // row 5, col 15

     reg start_in_5_15;
     wire start_out_5_15;

     reg [1:0] op_in_5_15;
     wire [1:0] op_out_5_15;

     wire r_5_15;

     reg data_in_5_15;
     wire data_out_5_15;

     reg pivot_in_5_15;
     wire pivot_out_5_15;

     always @(posedge clk) begin
         op_in_5_15 <= op_out_5_14;
         pivot_in_5_15 <= pivot_out_5_14;
         start_in_5_15 <= start_out_5_14;
     end

     always @(posedge clk) begin
         data_in_5_15 <= data_out_4_15;
     end
  
     processor_AB AB_5_15 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_15),
       .start_in   (start_in_5_15),
       .op_in      (op_in_5_15),
       .pivot_in   (pivot_in_5_15),
       .start_out  (start_out_5_15),
       .data_out   (data_out_5_15),
       .op_out     (op_out_5_15),
       .pivot_out  (pivot_out_5_15),
       .r          (r_5_15)
     );

  // row 5, col 16

     reg start_in_5_16;
     wire start_out_5_16;

     reg [1:0] op_in_5_16;
     wire [1:0] op_out_5_16;

     wire r_5_16;

     reg data_in_5_16;
     wire data_out_5_16;

     reg pivot_in_5_16;
     wire pivot_out_5_16;

     always @(posedge clk) begin
         op_in_5_16 <= op_out_5_15;
         pivot_in_5_16 <= pivot_out_5_15;
         start_in_5_16 <= start_out_5_15;
     end

     always @(posedge clk) begin
         data_in_5_16 <= data_out_4_16;
     end
  
     processor_AB AB_5_16 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_16),
       .start_in   (start_in_5_16),
       .op_in      (op_in_5_16),
       .pivot_in   (pivot_in_5_16),
       .start_out  (start_out_5_16),
       .data_out   (data_out_5_16),
       .op_out     (op_out_5_16),
       .pivot_out  (pivot_out_5_16),
       .r          (r_5_16)
     );

  // row 5, col 17

     reg start_in_5_17;
     wire start_out_5_17;

     reg [1:0] op_in_5_17;
     wire [1:0] op_out_5_17;

     wire r_5_17;

     reg data_in_5_17;
     wire data_out_5_17;

     reg pivot_in_5_17;
     wire pivot_out_5_17;

     always @(posedge clk) begin
         op_in_5_17 <= op_out_5_16;
         pivot_in_5_17 <= pivot_out_5_16;
         start_in_5_17 <= start_out_5_16;
     end

     always @(posedge clk) begin
         data_in_5_17 <= data_out_4_17;
     end
  
     processor_AB AB_5_17 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_17),
       .start_in   (start_in_5_17),
       .op_in      (op_in_5_17),
       .pivot_in   (pivot_in_5_17),
       .start_out  (start_out_5_17),
       .data_out   (data_out_5_17),
       .op_out     (op_out_5_17),
       .pivot_out  (pivot_out_5_17),
       .r          (r_5_17)
     );

  // row 5, col 18

     reg start_in_5_18;
     wire start_out_5_18;

     reg [1:0] op_in_5_18;
     wire [1:0] op_out_5_18;

     wire r_5_18;

     reg data_in_5_18;
     wire data_out_5_18;

     reg pivot_in_5_18;
     wire pivot_out_5_18;

     always @(posedge clk) begin
         op_in_5_18 <= op_out_5_17;
         pivot_in_5_18 <= pivot_out_5_17;
         start_in_5_18 <= start_out_5_17;
     end

     always @(posedge clk) begin
         data_in_5_18 <= data_out_4_18;
     end
  
     processor_AB AB_5_18 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_18),
       .start_in   (start_in_5_18),
       .op_in      (op_in_5_18),
       .pivot_in   (pivot_in_5_18),
       .start_out  (start_out_5_18),
       .data_out   (data_out_5_18),
       .op_out     (op_out_5_18),
       .pivot_out  (pivot_out_5_18),
       .r          (r_5_18)
     );

  // row 5, col 19

     reg start_in_5_19;
     wire start_out_5_19;

     reg [1:0] op_in_5_19;
     wire [1:0] op_out_5_19;

     wire r_5_19;

     reg data_in_5_19;
     wire data_out_5_19;

     reg pivot_in_5_19;
     wire pivot_out_5_19;

     always @(posedge clk) begin
         op_in_5_19 <= op_out_5_18;
         pivot_in_5_19 <= pivot_out_5_18;
         start_in_5_19 <= start_out_5_18;
     end

     always @(posedge clk) begin
         data_in_5_19 <= data_out_4_19;
     end
  
     processor_AB AB_5_19 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_19),
       .start_in   (start_in_5_19),
       .op_in      (op_in_5_19),
       .pivot_in   (pivot_in_5_19),
       .start_out  (start_out_5_19),
       .data_out   (data_out_5_19),
       .op_out     (op_out_5_19),
       .pivot_out  (pivot_out_5_19),
       .r          (r_5_19)
     );

  // row 5, col 20

     reg start_in_5_20;
     wire start_out_5_20;

     reg [1:0] op_in_5_20;
     wire [1:0] op_out_5_20;

     wire r_5_20;

     reg data_in_5_20;
     wire data_out_5_20;

     reg pivot_in_5_20;
     wire pivot_out_5_20;

     always @(posedge clk) begin
         op_in_5_20 <= op_out_5_19;
         pivot_in_5_20 <= pivot_out_5_19;
         start_in_5_20 <= start_out_5_19;
     end

     always @(posedge clk) begin
         data_in_5_20 <= data_out_4_20;
     end
  
     processor_AB AB_5_20 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_20),
       .start_in   (start_in_5_20),
       .op_in      (op_in_5_20),
       .pivot_in   (pivot_in_5_20),
       .start_out  (start_out_5_20),
       .data_out   (data_out_5_20),
       .op_out     (op_out_5_20),
       .pivot_out  (pivot_out_5_20),
       .r          (r_5_20)
     );

  // row 5, col 21

     reg start_in_5_21;
     wire start_out_5_21;

     reg [1:0] op_in_5_21;
     wire [1:0] op_out_5_21;

     wire r_5_21;

     reg data_in_5_21;
     wire data_out_5_21;

     reg pivot_in_5_21;
     wire pivot_out_5_21;

     always @(posedge clk) begin
         op_in_5_21 <= op_out_5_20;
         pivot_in_5_21 <= pivot_out_5_20;
         start_in_5_21 <= start_out_5_20;
     end

     always @(posedge clk) begin
         data_in_5_21 <= data_out_4_21;
     end
  
     processor_AB AB_5_21 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_21),
       .start_in   (start_in_5_21),
       .op_in      (op_in_5_21),
       .pivot_in   (pivot_in_5_21),
       .start_out  (start_out_5_21),
       .data_out   (data_out_5_21),
       .op_out     (op_out_5_21),
       .pivot_out  (pivot_out_5_21),
       .r          (r_5_21)
     );

  // row 5, col 22

     reg start_in_5_22;
     wire start_out_5_22;

     reg [1:0] op_in_5_22;
     wire [1:0] op_out_5_22;

     wire r_5_22;

     reg data_in_5_22;
     wire data_out_5_22;

     reg pivot_in_5_22;
     wire pivot_out_5_22;

     always @(posedge clk) begin
         op_in_5_22 <= op_out_5_21;
         pivot_in_5_22 <= pivot_out_5_21;
         start_in_5_22 <= start_out_5_21;
     end

     always @(posedge clk) begin
         data_in_5_22 <= data_out_4_22;
     end
  
     processor_AB AB_5_22 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_22),
       .start_in   (start_in_5_22),
       .op_in      (op_in_5_22),
       .pivot_in   (pivot_in_5_22),
       .start_out  (start_out_5_22),
       .data_out   (data_out_5_22),
       .op_out     (op_out_5_22),
       .pivot_out  (pivot_out_5_22),
       .r          (r_5_22)
     );

  // row 5, col 23

     reg start_in_5_23;
     wire start_out_5_23;

     reg [1:0] op_in_5_23;
     wire [1:0] op_out_5_23;

     wire r_5_23;

     reg data_in_5_23;
     wire data_out_5_23;

     reg pivot_in_5_23;
     wire pivot_out_5_23;

     always @(posedge clk) begin
         op_in_5_23 <= op_out_5_22;
         pivot_in_5_23 <= pivot_out_5_22;
         start_in_5_23 <= start_out_5_22;
     end

     always @(posedge clk) begin
         data_in_5_23 <= data_out_4_23;
     end
  
     processor_AB AB_5_23 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_23),
       .start_in   (start_in_5_23),
       .op_in      (op_in_5_23),
       .pivot_in   (pivot_in_5_23),
       .start_out  (start_out_5_23),
       .data_out   (data_out_5_23),
       .op_out     (op_out_5_23),
       .pivot_out  (pivot_out_5_23),
       .r          (r_5_23)
     );

  // row 5, col 24

     reg start_in_5_24;
     wire start_out_5_24;

     reg [1:0] op_in_5_24;
     wire [1:0] op_out_5_24;

     wire r_5_24;

     reg data_in_5_24;
     wire data_out_5_24;

     reg pivot_in_5_24;
     wire pivot_out_5_24;

     always @(posedge clk) begin
         op_in_5_24 <= op_out_5_23;
         pivot_in_5_24 <= pivot_out_5_23;
         start_in_5_24 <= start_out_5_23;
     end

     always @(posedge clk) begin
         data_in_5_24 <= data_out_4_24;
     end
  
     processor_AB AB_5_24 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_24),
       .start_in   (start_in_5_24),
       .op_in      (op_in_5_24),
       .pivot_in   (pivot_in_5_24),
       .start_out  (start_out_5_24),
       .data_out   (data_out_5_24),
       .op_out     (op_out_5_24),
       .pivot_out  (pivot_out_5_24),
       .r          (r_5_24)
     );

  // row 5, col 25

     reg start_in_5_25;
     wire start_out_5_25;

     reg [1:0] op_in_5_25;
     wire [1:0] op_out_5_25;

     wire r_5_25;

     reg data_in_5_25;
     wire data_out_5_25;

     reg pivot_in_5_25;
     wire pivot_out_5_25;

     always @(posedge clk) begin
         op_in_5_25 <= op_out_5_24;
         pivot_in_5_25 <= pivot_out_5_24;
         start_in_5_25 <= start_out_5_24;
     end

     always @(posedge clk) begin
         data_in_5_25 <= data_out_4_25;
     end
  
     processor_AB AB_5_25 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_25),
       .start_in   (start_in_5_25),
       .op_in      (op_in_5_25),
       .pivot_in   (pivot_in_5_25),
       .start_out  (start_out_5_25),
       .data_out   (data_out_5_25),
       .op_out     (op_out_5_25),
       .pivot_out  (pivot_out_5_25),
       .r          (r_5_25)
     );

  // row 5, col 26

     reg start_in_5_26;
     wire start_out_5_26;

     reg [1:0] op_in_5_26;
     wire [1:0] op_out_5_26;

     wire r_5_26;

     reg data_in_5_26;
     wire data_out_5_26;

     reg pivot_in_5_26;
     wire pivot_out_5_26;

     always @(posedge clk) begin
         op_in_5_26 <= op_out_5_25;
         pivot_in_5_26 <= pivot_out_5_25;
         start_in_5_26 <= start_out_5_25;
     end

     always @(posedge clk) begin
         data_in_5_26 <= data_out_4_26;
     end
  
     processor_AB AB_5_26 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_26),
       .start_in   (start_in_5_26),
       .op_in      (op_in_5_26),
       .pivot_in   (pivot_in_5_26),
       .start_out  (start_out_5_26),
       .data_out   (data_out_5_26),
       .op_out     (op_out_5_26),
       .pivot_out  (pivot_out_5_26),
       .r          (r_5_26)
     );

  // row 5, col 27

     reg start_in_5_27;
     wire start_out_5_27;

     reg [1:0] op_in_5_27;
     wire [1:0] op_out_5_27;

     wire r_5_27;

     reg data_in_5_27;
     wire data_out_5_27;

     reg pivot_in_5_27;
     wire pivot_out_5_27;

     always @(posedge clk) begin
         op_in_5_27 <= op_out_5_26;
         pivot_in_5_27 <= pivot_out_5_26;
         start_in_5_27 <= start_out_5_26;
     end

     always @(posedge clk) begin
         data_in_5_27 <= data_out_4_27;
     end
  
     processor_AB AB_5_27 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_27),
       .start_in   (start_in_5_27),
       .op_in      (op_in_5_27),
       .pivot_in   (pivot_in_5_27),
       .start_out  (start_out_5_27),
       .data_out   (data_out_5_27),
       .op_out     (op_out_5_27),
       .pivot_out  (pivot_out_5_27),
       .r          (r_5_27)
     );

  // row 5, col 28

     reg start_in_5_28;
     wire start_out_5_28;

     reg [1:0] op_in_5_28;
     wire [1:0] op_out_5_28;

     wire r_5_28;

     reg data_in_5_28;
     wire data_out_5_28;

     reg pivot_in_5_28;
     wire pivot_out_5_28;

     always @(posedge clk) begin
         op_in_5_28 <= op_out_5_27;
         pivot_in_5_28 <= pivot_out_5_27;
         start_in_5_28 <= start_out_5_27;
     end

     always @(posedge clk) begin
         data_in_5_28 <= data_out_4_28;
     end
  
     processor_AB AB_5_28 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_28),
       .start_in   (start_in_5_28),
       .op_in      (op_in_5_28),
       .pivot_in   (pivot_in_5_28),
       .start_out  (start_out_5_28),
       .data_out   (data_out_5_28),
       .op_out     (op_out_5_28),
       .pivot_out  (pivot_out_5_28),
       .r          (r_5_28)
     );

  // row 5, col 29

     reg start_in_5_29;
     wire start_out_5_29;

     reg [1:0] op_in_5_29;
     wire [1:0] op_out_5_29;

     wire r_5_29;

     reg data_in_5_29;
     wire data_out_5_29;

     reg pivot_in_5_29;
     wire pivot_out_5_29;

     always @(posedge clk) begin
         op_in_5_29 <= op_out_5_28;
         pivot_in_5_29 <= pivot_out_5_28;
         start_in_5_29 <= start_out_5_28;
     end

     always @(posedge clk) begin
         data_in_5_29 <= data_out_4_29;
     end
  
     processor_AB AB_5_29 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_29),
       .start_in   (start_in_5_29),
       .op_in      (op_in_5_29),
       .pivot_in   (pivot_in_5_29),
       .start_out  (start_out_5_29),
       .data_out   (data_out_5_29),
       .op_out     (op_out_5_29),
       .pivot_out  (pivot_out_5_29),
       .r          (r_5_29)
     );

  // row 5, col 30

     reg start_in_5_30;
     wire start_out_5_30;

     reg [1:0] op_in_5_30;
     wire [1:0] op_out_5_30;

     wire r_5_30;

     reg data_in_5_30;
     wire data_out_5_30;

     reg pivot_in_5_30;
     wire pivot_out_5_30;

     always @(posedge clk) begin
         op_in_5_30 <= op_out_5_29;
         pivot_in_5_30 <= pivot_out_5_29;
         start_in_5_30 <= start_out_5_29;
     end

     always @(posedge clk) begin
         data_in_5_30 <= data_out_4_30;
     end
  
     processor_AB AB_5_30 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_30),
       .start_in   (start_in_5_30),
       .op_in      (op_in_5_30),
       .pivot_in   (pivot_in_5_30),
       .start_out  (start_out_5_30),
       .data_out   (data_out_5_30),
       .op_out     (op_out_5_30),
       .pivot_out  (pivot_out_5_30),
       .r          (r_5_30)
     );

  // row 5, col 31

     reg start_in_5_31;
     wire start_out_5_31;

     reg [1:0] op_in_5_31;
     wire [1:0] op_out_5_31;

     wire r_5_31;

     reg data_in_5_31;
     wire data_out_5_31;

     reg pivot_in_5_31;
     wire pivot_out_5_31;

     always @(posedge clk) begin
         op_in_5_31 <= op_out_5_30;
         pivot_in_5_31 <= pivot_out_5_30;
         start_in_5_31 <= start_out_5_30;
     end

     always @(posedge clk) begin
         data_in_5_31 <= data_out_4_31;
     end
  
     processor_AB AB_5_31 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_31),
       .start_in   (start_in_5_31),
       .op_in      (op_in_5_31),
       .pivot_in   (pivot_in_5_31),
       .start_out  (start_out_5_31),
       .data_out   (data_out_5_31),
       .op_out     (op_out_5_31),
       .pivot_out  (pivot_out_5_31),
       .r          (r_5_31)
     );

  // row 5, col 32

     reg start_in_5_32;
     wire start_out_5_32;

     reg [1:0] op_in_5_32;
     wire [1:0] op_out_5_32;

     wire r_5_32;

     reg data_in_5_32;
     wire data_out_5_32;

     reg pivot_in_5_32;
     wire pivot_out_5_32;

     always @(posedge clk) begin
         op_in_5_32 <= op_out_5_31;
         pivot_in_5_32 <= pivot_out_5_31;
         start_in_5_32 <= start_out_5_31;
     end

     always @(posedge clk) begin
         data_in_5_32 <= data_out_4_32;
     end
  
     processor_AB AB_5_32 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_32),
       .start_in   (start_in_5_32),
       .op_in      (op_in_5_32),
       .pivot_in   (pivot_in_5_32),
       .start_out  (start_out_5_32),
       .data_out   (data_out_5_32),
       .op_out     (op_out_5_32),
       .pivot_out  (pivot_out_5_32),
       .r          (r_5_32)
     );

  // row 5, col 33

     reg start_in_5_33;
     wire start_out_5_33;

     reg [1:0] op_in_5_33;
     wire [1:0] op_out_5_33;

     wire r_5_33;

     reg data_in_5_33;
     wire data_out_5_33;

     reg pivot_in_5_33;
     wire pivot_out_5_33;

     always @(posedge clk) begin
         op_in_5_33 <= op_out_5_32;
         pivot_in_5_33 <= pivot_out_5_32;
         start_in_5_33 <= start_out_5_32;
     end

     always @(posedge clk) begin
         data_in_5_33 <= data_out_4_33;
     end
  
     processor_AB AB_5_33 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_33),
       .start_in   (start_in_5_33),
       .op_in      (op_in_5_33),
       .pivot_in   (pivot_in_5_33),
       .start_out  (start_out_5_33),
       .data_out   (data_out_5_33),
       .op_out     (op_out_5_33),
       .pivot_out  (pivot_out_5_33),
       .r          (r_5_33)
     );

  // row 5, col 34

     reg start_in_5_34;
     wire start_out_5_34;

     reg [1:0] op_in_5_34;
     wire [1:0] op_out_5_34;

     wire r_5_34;

     reg data_in_5_34;
     wire data_out_5_34;

     reg pivot_in_5_34;
     wire pivot_out_5_34;

     always @(posedge clk) begin
         op_in_5_34 <= op_out_5_33;
         pivot_in_5_34 <= pivot_out_5_33;
         start_in_5_34 <= start_out_5_33;
     end

     always @(posedge clk) begin
         data_in_5_34 <= data_out_4_34;
     end
  
     processor_AB AB_5_34 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_34),
       .start_in   (start_in_5_34),
       .op_in      (op_in_5_34),
       .pivot_in   (pivot_in_5_34),
       .start_out  (start_out_5_34),
       .data_out   (data_out_5_34),
       .op_out     (op_out_5_34),
       .pivot_out  (pivot_out_5_34),
       .r          (r_5_34)
     );

  // row 5, col 35

     reg start_in_5_35;
     wire start_out_5_35;

     reg [1:0] op_in_5_35;
     wire [1:0] op_out_5_35;

     wire r_5_35;

     reg data_in_5_35;
     wire data_out_5_35;

     reg pivot_in_5_35;
     wire pivot_out_5_35;

     always @(posedge clk) begin
         op_in_5_35 <= op_out_5_34;
         pivot_in_5_35 <= pivot_out_5_34;
         start_in_5_35 <= start_out_5_34;
     end

     always @(posedge clk) begin
         data_in_5_35 <= data_out_4_35;
     end
  
     processor_AB AB_5_35 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_35),
       .start_in   (start_in_5_35),
       .op_in      (op_in_5_35),
       .pivot_in   (pivot_in_5_35),
       .start_out  (start_out_5_35),
       .data_out   (data_out_5_35),
       .op_out     (op_out_5_35),
       .pivot_out  (pivot_out_5_35),
       .r          (r_5_35)
     );

  // row 5, col 36

     reg start_in_5_36;
     wire start_out_5_36;

     reg [1:0] op_in_5_36;
     wire [1:0] op_out_5_36;

     wire r_5_36;

     reg data_in_5_36;
     wire data_out_5_36;

     reg pivot_in_5_36;
     wire pivot_out_5_36;

     always @(posedge clk) begin
         op_in_5_36 <= op_out_5_35;
         pivot_in_5_36 <= pivot_out_5_35;
         start_in_5_36 <= start_out_5_35;
     end

     always @(posedge clk) begin
         data_in_5_36 <= data_out_4_36;
     end
  
     processor_AB AB_5_36 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_36),
       .start_in   (start_in_5_36),
       .op_in      (op_in_5_36),
       .pivot_in   (pivot_in_5_36),
       .start_out  (start_out_5_36),
       .data_out   (data_out_5_36),
       .op_out     (op_out_5_36),
       .pivot_out  (pivot_out_5_36),
       .r          (r_5_36)
     );

  // row 5, col 37

     reg start_in_5_37;
     wire start_out_5_37;

     reg [1:0] op_in_5_37;
     wire [1:0] op_out_5_37;

     wire r_5_37;

     reg data_in_5_37;
     wire data_out_5_37;

     reg pivot_in_5_37;
     wire pivot_out_5_37;

     always @(posedge clk) begin
         op_in_5_37 <= op_out_5_36;
         pivot_in_5_37 <= pivot_out_5_36;
         start_in_5_37 <= start_out_5_36;
     end

     always @(posedge clk) begin
         data_in_5_37 <= data_out_4_37;
     end
  
     processor_AB AB_5_37 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_37),
       .start_in   (start_in_5_37),
       .op_in      (op_in_5_37),
       .pivot_in   (pivot_in_5_37),
       .start_out  (start_out_5_37),
       .data_out   (data_out_5_37),
       .op_out     (op_out_5_37),
       .pivot_out  (pivot_out_5_37),
       .r          (r_5_37)
     );

  // row 5, col 38

     reg start_in_5_38;
     wire start_out_5_38;

     reg [1:0] op_in_5_38;
     wire [1:0] op_out_5_38;

     wire r_5_38;

     reg data_in_5_38;
     wire data_out_5_38;

     reg pivot_in_5_38;
     wire pivot_out_5_38;

     always @(posedge clk) begin
         op_in_5_38 <= op_out_5_37;
         pivot_in_5_38 <= pivot_out_5_37;
         start_in_5_38 <= start_out_5_37;
     end

     always @(posedge clk) begin
         data_in_5_38 <= data_out_4_38;
     end
  
     processor_AB AB_5_38 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_38),
       .start_in   (start_in_5_38),
       .op_in      (op_in_5_38),
       .pivot_in   (pivot_in_5_38),
       .start_out  (start_out_5_38),
       .data_out   (data_out_5_38),
       .op_out     (op_out_5_38),
       .pivot_out  (pivot_out_5_38),
       .r          (r_5_38)
     );

  // row 5, col 39

     reg start_in_5_39;
     wire start_out_5_39;

     reg [1:0] op_in_5_39;
     wire [1:0] op_out_5_39;

     wire r_5_39;

     reg data_in_5_39;
     wire data_out_5_39;

     reg pivot_in_5_39;
     wire pivot_out_5_39;

     always @(posedge clk) begin
         op_in_5_39 <= op_out_5_38;
         pivot_in_5_39 <= pivot_out_5_38;
         start_in_5_39 <= start_out_5_38;
     end

     always @(posedge clk) begin
         data_in_5_39 <= data_out_4_39;
     end
  
     processor_AB AB_5_39 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_39),
       .start_in   (start_in_5_39),
       .op_in      (op_in_5_39),
       .pivot_in   (pivot_in_5_39),
       .start_out  (start_out_5_39),
       .data_out   (data_out_5_39),
       .op_out     (op_out_5_39),
       .pivot_out  (pivot_out_5_39),
       .r          (r_5_39)
     );

  // row 5, col 40

     reg start_in_5_40;
     wire start_out_5_40;

     reg [1:0] op_in_5_40;
     wire [1:0] op_out_5_40;

     wire r_5_40;

     reg data_in_5_40;
     wire data_out_5_40;

     reg pivot_in_5_40;
     wire pivot_out_5_40;

     always @(posedge clk) begin
         op_in_5_40 <= op_out_5_39;
         pivot_in_5_40 <= pivot_out_5_39;
         start_in_5_40 <= start_out_5_39;
     end

     always @(posedge clk) begin
         data_in_5_40 <= data_out_4_40;
     end
  
     processor_AB AB_5_40 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_40),
       .start_in   (start_in_5_40),
       .op_in      (op_in_5_40),
       .pivot_in   (pivot_in_5_40),
       .start_out  (start_out_5_40),
       .data_out   (data_out_5_40),
       .op_out     (op_out_5_40),
       .pivot_out  (pivot_out_5_40),
       .r          (r_5_40)
     );

  // row 5, col 41

     reg start_in_5_41;
     wire start_out_5_41;

     reg [1:0] op_in_5_41;
     wire [1:0] op_out_5_41;

     wire r_5_41;

     reg data_in_5_41;
     wire data_out_5_41;

     reg pivot_in_5_41;
     wire pivot_out_5_41;

     always @(posedge clk) begin
         op_in_5_41 <= op_out_5_40;
         pivot_in_5_41 <= pivot_out_5_40;
         start_in_5_41 <= start_out_5_40;
     end

     always @(posedge clk) begin
         data_in_5_41 <= data_out_4_41;
     end
  
     processor_AB AB_5_41 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_41),
       .start_in   (start_in_5_41),
       .op_in      (op_in_5_41),
       .pivot_in   (pivot_in_5_41),
       .start_out  (start_out_5_41),
       .data_out   (data_out_5_41),
       .op_out     (op_out_5_41),
       .pivot_out  (pivot_out_5_41),
       .r          (r_5_41)
     );

  // row 5, col 42

     reg start_in_5_42;
     wire start_out_5_42;

     reg [1:0] op_in_5_42;
     wire [1:0] op_out_5_42;

     wire r_5_42;

     reg data_in_5_42;
     wire data_out_5_42;

     reg pivot_in_5_42;
     wire pivot_out_5_42;

     always @(posedge clk) begin
         op_in_5_42 <= op_out_5_41;
         pivot_in_5_42 <= pivot_out_5_41;
         start_in_5_42 <= start_out_5_41;
     end

     always @(posedge clk) begin
         data_in_5_42 <= data_out_4_42;
     end
  
     processor_AB AB_5_42 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_42),
       .start_in   (start_in_5_42),
       .op_in      (op_in_5_42),
       .pivot_in   (pivot_in_5_42),
       .start_out  (start_out_5_42),
       .data_out   (data_out_5_42),
       .op_out     (op_out_5_42),
       .pivot_out  (pivot_out_5_42),
       .r          (r_5_42)
     );

  // row 5, col 43

     reg start_in_5_43;
     wire start_out_5_43;

     reg [1:0] op_in_5_43;
     wire [1:0] op_out_5_43;

     wire r_5_43;

     reg data_in_5_43;
     wire data_out_5_43;

     reg pivot_in_5_43;
     wire pivot_out_5_43;

     always @(posedge clk) begin
         op_in_5_43 <= op_out_5_42;
         pivot_in_5_43 <= pivot_out_5_42;
         start_in_5_43 <= start_out_5_42;
     end

     always @(posedge clk) begin
         data_in_5_43 <= data_out_4_43;
     end
  
     processor_AB AB_5_43 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_43),
       .start_in   (start_in_5_43),
       .op_in      (op_in_5_43),
       .pivot_in   (pivot_in_5_43),
       .start_out  (start_out_5_43),
       .data_out   (data_out_5_43),
       .op_out     (op_out_5_43),
       .pivot_out  (pivot_out_5_43),
       .r          (r_5_43)
     );

  // row 5, col 44

     reg start_in_5_44;
     wire start_out_5_44;

     reg [1:0] op_in_5_44;
     wire [1:0] op_out_5_44;

     wire r_5_44;

     reg data_in_5_44;
     wire data_out_5_44;

     reg pivot_in_5_44;
     wire pivot_out_5_44;

     always @(posedge clk) begin
         op_in_5_44 <= op_out_5_43;
         pivot_in_5_44 <= pivot_out_5_43;
         start_in_5_44 <= start_out_5_43;
     end

     always @(posedge clk) begin
         data_in_5_44 <= data_out_4_44;
     end
  
     processor_AB AB_5_44 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_44),
       .start_in   (start_in_5_44),
       .op_in      (op_in_5_44),
       .pivot_in   (pivot_in_5_44),
       .start_out  (start_out_5_44),
       .data_out   (data_out_5_44),
       .op_out     (op_out_5_44),
       .pivot_out  (pivot_out_5_44),
       .r          (r_5_44)
     );

  // row 5, col 45

     reg start_in_5_45;
     wire start_out_5_45;

     reg [1:0] op_in_5_45;
     wire [1:0] op_out_5_45;

     wire r_5_45;

     reg data_in_5_45;
     wire data_out_5_45;

     reg pivot_in_5_45;
     wire pivot_out_5_45;

     always @(posedge clk) begin
         op_in_5_45 <= op_out_5_44;
         pivot_in_5_45 <= pivot_out_5_44;
         start_in_5_45 <= start_out_5_44;
     end

     always @(posedge clk) begin
         data_in_5_45 <= data_out_4_45;
     end
  
     processor_AB AB_5_45 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_45),
       .start_in   (start_in_5_45),
       .op_in      (op_in_5_45),
       .pivot_in   (pivot_in_5_45),
       .start_out  (start_out_5_45),
       .data_out   (data_out_5_45),
       .op_out     (op_out_5_45),
       .pivot_out  (pivot_out_5_45),
       .r          (r_5_45)
     );

  // row 5, col 46

     reg start_in_5_46;
     wire start_out_5_46;

     reg [1:0] op_in_5_46;
     wire [1:0] op_out_5_46;

     wire r_5_46;

     reg data_in_5_46;
     wire data_out_5_46;

     reg pivot_in_5_46;
     wire pivot_out_5_46;

     always @(posedge clk) begin
         op_in_5_46 <= op_out_5_45;
         pivot_in_5_46 <= pivot_out_5_45;
         start_in_5_46 <= start_out_5_45;
     end

     always @(posedge clk) begin
         data_in_5_46 <= data_out_4_46;
     end
  
     processor_AB AB_5_46 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_46),
       .start_in   (start_in_5_46),
       .op_in      (op_in_5_46),
       .pivot_in   (pivot_in_5_46),
       .start_out  (start_out_5_46),
       .data_out   (data_out_5_46),
       .op_out     (op_out_5_46),
       .pivot_out  (pivot_out_5_46),
       .r          (r_5_46)
     );

  // row 5, col 47

     reg start_in_5_47;
     wire start_out_5_47;

     reg [1:0] op_in_5_47;
     wire [1:0] op_out_5_47;

     wire r_5_47;

     reg data_in_5_47;
     wire data_out_5_47;

     reg pivot_in_5_47;
     wire pivot_out_5_47;

     always @(posedge clk) begin
         op_in_5_47 <= op_out_5_46;
         pivot_in_5_47 <= pivot_out_5_46;
         start_in_5_47 <= start_out_5_46;
     end

     always @(posedge clk) begin
         data_in_5_47 <= data_out_4_47;
     end
  
     processor_AB AB_5_47 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_47),
       .start_in   (start_in_5_47),
       .op_in      (op_in_5_47),
       .pivot_in   (pivot_in_5_47),
       .start_out  (start_out_5_47),
       .data_out   (data_out_5_47),
       .op_out     (op_out_5_47),
       .pivot_out  (pivot_out_5_47),
       .r          (r_5_47)
     );

  // row 5, col 48

     reg start_in_5_48;
     wire start_out_5_48;

     reg [1:0] op_in_5_48;
     wire [1:0] op_out_5_48;

     wire r_5_48;

     reg data_in_5_48;
     wire data_out_5_48;

     reg pivot_in_5_48;
     wire pivot_out_5_48;

     always @(posedge clk) begin
         op_in_5_48 <= op_out_5_47;
         pivot_in_5_48 <= pivot_out_5_47;
         start_in_5_48 <= start_out_5_47;
     end

     always @(posedge clk) begin
         data_in_5_48 <= data_out_4_48;
     end
  
     processor_AB AB_5_48 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_48),
       .start_in   (start_in_5_48),
       .op_in      (op_in_5_48),
       .pivot_in   (pivot_in_5_48),
       .start_out  (start_out_5_48),
       .data_out   (data_out_5_48),
       .op_out     (op_out_5_48),
       .pivot_out  (pivot_out_5_48),
       .r          (r_5_48)
     );

  // row 5, col 49

     reg start_in_5_49;
     wire start_out_5_49;

     reg [1:0] op_in_5_49;
     wire [1:0] op_out_5_49;

     wire r_5_49;

     reg data_in_5_49;
     wire data_out_5_49;

     reg pivot_in_5_49;
     wire pivot_out_5_49;

     always @(posedge clk) begin
         op_in_5_49 <= op_out_5_48;
         pivot_in_5_49 <= pivot_out_5_48;
         start_in_5_49 <= start_out_5_48;
     end

     always @(posedge clk) begin
         data_in_5_49 <= data_out_4_49;
     end
  
     processor_AB AB_5_49 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_49),
       .start_in   (start_in_5_49),
       .op_in      (op_in_5_49),
       .pivot_in   (pivot_in_5_49),
       .start_out  (start_out_5_49),
       .data_out   (data_out_5_49),
       .op_out     (op_out_5_49),
       .pivot_out  (pivot_out_5_49),
       .r          (r_5_49)
     );

  // row 5, col 50

     reg start_in_5_50;
     wire start_out_5_50;

     reg [1:0] op_in_5_50;
     wire [1:0] op_out_5_50;

     wire r_5_50;

     reg data_in_5_50;
     wire data_out_5_50;

     reg pivot_in_5_50;
     wire pivot_out_5_50;

     always @(posedge clk) begin
         op_in_5_50 <= op_out_5_49;
         pivot_in_5_50 <= pivot_out_5_49;
         start_in_5_50 <= start_out_5_49;
     end

     always @(posedge clk) begin
         data_in_5_50 <= data_out_4_50;
     end
  
     processor_AB AB_5_50 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_50),
       .start_in   (start_in_5_50),
       .op_in      (op_in_5_50),
       .pivot_in   (pivot_in_5_50),
       .start_out  (start_out_5_50),
       .data_out   (data_out_5_50),
       .op_out     (op_out_5_50),
       .pivot_out  (pivot_out_5_50),
       .r          (r_5_50)
     );

  // row 5, col 51

     reg start_in_5_51;
     wire start_out_5_51;

     reg [1:0] op_in_5_51;
     wire [1:0] op_out_5_51;

     wire r_5_51;

     reg data_in_5_51;
     wire data_out_5_51;

     reg pivot_in_5_51;
     wire pivot_out_5_51;

     always @(posedge clk) begin
         op_in_5_51 <= op_out_5_50;
         pivot_in_5_51 <= pivot_out_5_50;
         start_in_5_51 <= start_out_5_50;
     end

     always @(posedge clk) begin
         data_in_5_51 <= data_out_4_51;
     end
  
     processor_AB AB_5_51 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_51),
       .start_in   (start_in_5_51),
       .op_in      (op_in_5_51),
       .pivot_in   (pivot_in_5_51),
       .start_out  (start_out_5_51),
       .data_out   (data_out_5_51),
       .op_out     (op_out_5_51),
       .pivot_out  (pivot_out_5_51),
       .r          (r_5_51)
     );

  // row 5, col 52

     reg start_in_5_52;
     wire start_out_5_52;

     reg [1:0] op_in_5_52;
     wire [1:0] op_out_5_52;

     wire r_5_52;

     reg data_in_5_52;
     wire data_out_5_52;

     reg pivot_in_5_52;
     wire pivot_out_5_52;

     always @(posedge clk) begin
         op_in_5_52 <= op_out_5_51;
         pivot_in_5_52 <= pivot_out_5_51;
         start_in_5_52 <= start_out_5_51;
     end

     always @(posedge clk) begin
         data_in_5_52 <= data_out_4_52;
     end
  
     processor_AB AB_5_52 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_52),
       .start_in   (start_in_5_52),
       .op_in      (op_in_5_52),
       .pivot_in   (pivot_in_5_52),
       .start_out  (start_out_5_52),
       .data_out   (data_out_5_52),
       .op_out     (op_out_5_52),
       .pivot_out  (pivot_out_5_52),
       .r          (r_5_52)
     );

  // row 5, col 53

     reg start_in_5_53;
     wire start_out_5_53;

     reg [1:0] op_in_5_53;
     wire [1:0] op_out_5_53;

     wire r_5_53;

     reg data_in_5_53;
     wire data_out_5_53;

     reg pivot_in_5_53;
     wire pivot_out_5_53;

     always @(posedge clk) begin
         op_in_5_53 <= op_out_5_52;
         pivot_in_5_53 <= pivot_out_5_52;
         start_in_5_53 <= start_out_5_52;
     end

     always @(posedge clk) begin
         data_in_5_53 <= data_out_4_53;
     end
  
     processor_AB AB_5_53 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_53),
       .start_in   (start_in_5_53),
       .op_in      (op_in_5_53),
       .pivot_in   (pivot_in_5_53),
       .start_out  (start_out_5_53),
       .data_out   (data_out_5_53),
       .op_out     (op_out_5_53),
       .pivot_out  (pivot_out_5_53),
       .r          (r_5_53)
     );

  // row 5, col 54

     reg start_in_5_54;
     wire start_out_5_54;

     reg [1:0] op_in_5_54;
     wire [1:0] op_out_5_54;

     wire r_5_54;

     reg data_in_5_54;
     wire data_out_5_54;

     reg pivot_in_5_54;
     wire pivot_out_5_54;

     always @(posedge clk) begin
         op_in_5_54 <= op_out_5_53;
         pivot_in_5_54 <= pivot_out_5_53;
         start_in_5_54 <= start_out_5_53;
     end

     always @(posedge clk) begin
         data_in_5_54 <= data_out_4_54;
     end
  
     processor_AB AB_5_54 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_54),
       .start_in   (start_in_5_54),
       .op_in      (op_in_5_54),
       .pivot_in   (pivot_in_5_54),
       .start_out  (start_out_5_54),
       .data_out   (data_out_5_54),
       .op_out     (op_out_5_54),
       .pivot_out  (pivot_out_5_54),
       .r          (r_5_54)
     );

  // row 5, col 55

     reg start_in_5_55;
     wire start_out_5_55;

     reg [1:0] op_in_5_55;
     wire [1:0] op_out_5_55;

     wire r_5_55;

     reg data_in_5_55;
     wire data_out_5_55;

     reg pivot_in_5_55;
     wire pivot_out_5_55;

     always @(posedge clk) begin
         op_in_5_55 <= op_out_5_54;
         pivot_in_5_55 <= pivot_out_5_54;
         start_in_5_55 <= start_out_5_54;
     end

     always @(posedge clk) begin
         data_in_5_55 <= data_out_4_55;
     end
  
     processor_AB AB_5_55 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_55),
       .start_in   (start_in_5_55),
       .op_in      (op_in_5_55),
       .pivot_in   (pivot_in_5_55),
       .start_out  (start_out_5_55),
       .data_out   (data_out_5_55),
       .op_out     (op_out_5_55),
       .pivot_out  (pivot_out_5_55),
       .r          (r_5_55)
     );

  // row 5, col 56

     reg start_in_5_56;
     wire start_out_5_56;

     reg [1:0] op_in_5_56;
     wire [1:0] op_out_5_56;

     wire r_5_56;

     reg data_in_5_56;
     wire data_out_5_56;

     reg pivot_in_5_56;
     wire pivot_out_5_56;

     always @(posedge clk) begin
         op_in_5_56 <= op_out_5_55;
         pivot_in_5_56 <= pivot_out_5_55;
         start_in_5_56 <= start_out_5_55;
     end

     always @(posedge clk) begin
         data_in_5_56 <= data_out_4_56;
     end
  
     processor_AB AB_5_56 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_56),
       .start_in   (start_in_5_56),
       .op_in      (op_in_5_56),
       .pivot_in   (pivot_in_5_56),
       .start_out  (start_out_5_56),
       .data_out   (data_out_5_56),
       .op_out     (op_out_5_56),
       .pivot_out  (pivot_out_5_56),
       .r          (r_5_56)
     );

  // row 5, col 57

     reg start_in_5_57;
     wire start_out_5_57;

     reg [1:0] op_in_5_57;
     wire [1:0] op_out_5_57;

     wire r_5_57;

     reg data_in_5_57;
     wire data_out_5_57;

     reg pivot_in_5_57;
     wire pivot_out_5_57;

     always @(posedge clk) begin
         op_in_5_57 <= op_out_5_56;
         pivot_in_5_57 <= pivot_out_5_56;
         start_in_5_57 <= start_out_5_56;
     end

     always @(posedge clk) begin
         data_in_5_57 <= data_out_4_57;
     end
  
     processor_AB AB_5_57 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_57),
       .start_in   (start_in_5_57),
       .op_in      (op_in_5_57),
       .pivot_in   (pivot_in_5_57),
       .start_out  (start_out_5_57),
       .data_out   (data_out_5_57),
       .op_out     (op_out_5_57),
       .pivot_out  (pivot_out_5_57),
       .r          (r_5_57)
     );

  // row 5, col 58

     reg start_in_5_58;
     wire start_out_5_58;

     reg [1:0] op_in_5_58;
     wire [1:0] op_out_5_58;

     wire r_5_58;

     reg data_in_5_58;
     wire data_out_5_58;

     reg pivot_in_5_58;
     wire pivot_out_5_58;

     always @(posedge clk) begin
         op_in_5_58 <= op_out_5_57;
         pivot_in_5_58 <= pivot_out_5_57;
         start_in_5_58 <= start_out_5_57;
     end

     always @(posedge clk) begin
         data_in_5_58 <= data_out_4_58;
     end
  
     processor_AB AB_5_58 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_58),
       .start_in   (start_in_5_58),
       .op_in      (op_in_5_58),
       .pivot_in   (pivot_in_5_58),
       .start_out  (start_out_5_58),
       .data_out   (data_out_5_58),
       .op_out     (op_out_5_58),
       .pivot_out  (pivot_out_5_58),
       .r          (r_5_58)
     );

  // row 5, col 59

     reg start_in_5_59;
     wire start_out_5_59;

     reg [1:0] op_in_5_59;
     wire [1:0] op_out_5_59;

     wire r_5_59;

     reg data_in_5_59;
     wire data_out_5_59;

     reg pivot_in_5_59;
     wire pivot_out_5_59;

     always @(posedge clk) begin
         op_in_5_59 <= op_out_5_58;
         pivot_in_5_59 <= pivot_out_5_58;
         start_in_5_59 <= start_out_5_58;
     end

     always @(posedge clk) begin
         data_in_5_59 <= data_out_4_59;
     end
  
     processor_AB AB_5_59 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_59),
       .start_in   (start_in_5_59),
       .op_in      (op_in_5_59),
       .pivot_in   (pivot_in_5_59),
       .start_out  (start_out_5_59),
       .data_out   (data_out_5_59),
       .op_out     (op_out_5_59),
       .pivot_out  (pivot_out_5_59),
       .r          (r_5_59)
     );

  // row 5, col 60

     reg start_in_5_60;
     wire start_out_5_60;

     reg [1:0] op_in_5_60;
     wire [1:0] op_out_5_60;

     wire r_5_60;

     reg data_in_5_60;
     wire data_out_5_60;

     reg pivot_in_5_60;
     wire pivot_out_5_60;

     always @(posedge clk) begin
         op_in_5_60 <= op_out_5_59;
         pivot_in_5_60 <= pivot_out_5_59;
         start_in_5_60 <= start_out_5_59;
     end

     always @(posedge clk) begin
         data_in_5_60 <= data_out_4_60;
     end
  
     processor_AB AB_5_60 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_60),
       .start_in   (start_in_5_60),
       .op_in      (op_in_5_60),
       .pivot_in   (pivot_in_5_60),
       .start_out  (start_out_5_60),
       .data_out   (data_out_5_60),
       .op_out     (op_out_5_60),
       .pivot_out  (pivot_out_5_60),
       .r          (r_5_60)
     );

  // row 5, col 61

     reg start_in_5_61;
     wire start_out_5_61;

     reg [1:0] op_in_5_61;
     wire [1:0] op_out_5_61;

     wire r_5_61;

     reg data_in_5_61;
     wire data_out_5_61;

     reg pivot_in_5_61;
     wire pivot_out_5_61;

     always @(posedge clk) begin
         op_in_5_61 <= op_out_5_60;
         pivot_in_5_61 <= pivot_out_5_60;
         start_in_5_61 <= start_out_5_60;
     end

     always @(posedge clk) begin
         data_in_5_61 <= data_out_4_61;
     end
  
     processor_AB AB_5_61 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_61),
       .start_in   (start_in_5_61),
       .op_in      (op_in_5_61),
       .pivot_in   (pivot_in_5_61),
       .start_out  (start_out_5_61),
       .data_out   (data_out_5_61),
       .op_out     (op_out_5_61),
       .pivot_out  (pivot_out_5_61),
       .r          (r_5_61)
     );

  // row 5, col 62

     reg start_in_5_62;
     wire start_out_5_62;

     reg [1:0] op_in_5_62;
     wire [1:0] op_out_5_62;

     wire r_5_62;

     reg data_in_5_62;
     wire data_out_5_62;

     reg pivot_in_5_62;
     wire pivot_out_5_62;

     always @(posedge clk) begin
         op_in_5_62 <= op_out_5_61;
         pivot_in_5_62 <= pivot_out_5_61;
         start_in_5_62 <= start_out_5_61;
     end

     always @(posedge clk) begin
         data_in_5_62 <= data_out_4_62;
     end
  
     processor_AB AB_5_62 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_62),
       .start_in   (start_in_5_62),
       .op_in      (op_in_5_62),
       .pivot_in   (pivot_in_5_62),
       .start_out  (start_out_5_62),
       .data_out   (data_out_5_62),
       .op_out     (op_out_5_62),
       .pivot_out  (pivot_out_5_62),
       .r          (r_5_62)
     );

  // row 5, col 63

     reg start_in_5_63;
     wire start_out_5_63;

     reg [1:0] op_in_5_63;
     wire [1:0] op_out_5_63;

     wire r_5_63;

     reg data_in_5_63;
     wire data_out_5_63;

     reg pivot_in_5_63;
     wire pivot_out_5_63;

     always @(posedge clk) begin
         op_in_5_63 <= op_out_5_62;
         pivot_in_5_63 <= pivot_out_5_62;
         start_in_5_63 <= start_out_5_62;
     end

     always @(posedge clk) begin
         data_in_5_63 <= data_out_4_63;
     end
  
     processor_AB AB_5_63 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_63),
       .start_in   (start_in_5_63),
       .op_in      (op_in_5_63),
       .pivot_in   (pivot_in_5_63),
       .start_out  (start_out_5_63),
       .data_out   (data_out_5_63),
       .op_out     (op_out_5_63),
       .pivot_out  (pivot_out_5_63),
       .r          (r_5_63)
     );

  // row 5, col 64

     reg start_in_5_64;
     wire start_out_5_64;

     reg [1:0] op_in_5_64;
     wire [1:0] op_out_5_64;

     wire r_5_64;

     reg data_in_5_64;
     wire data_out_5_64;

     reg pivot_in_5_64;
     wire pivot_out_5_64;

     always @(posedge clk) begin
         op_in_5_64 <= op_out_5_63;
         pivot_in_5_64 <= pivot_out_5_63;
         start_in_5_64 <= start_out_5_63;
     end

     always @(posedge clk) begin
         data_in_5_64 <= data_out_4_64;
     end
  
     processor_AB AB_5_64 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_64),
       .start_in   (start_in_5_64),
       .op_in      (op_in_5_64),
       .pivot_in   (pivot_in_5_64),
       .start_out  (start_out_5_64),
       .data_out   (data_out_5_64),
       .op_out     (op_out_5_64),
       .pivot_out  (pivot_out_5_64),
       .r          (r_5_64)
     );

  // row 5, col 65

     reg start_in_5_65;
     wire start_out_5_65;

     reg [1:0] op_in_5_65;
     wire [1:0] op_out_5_65;

     wire r_5_65;

     reg data_in_5_65;
     wire data_out_5_65;

     reg pivot_in_5_65;
     wire pivot_out_5_65;

     always @(posedge clk) begin
         op_in_5_65 <= op_out_5_64;
         pivot_in_5_65 <= pivot_out_5_64;
         start_in_5_65 <= start_out_5_64;
     end

     always @(posedge clk) begin
         data_in_5_65 <= data_out_4_65;
     end
  
     processor_AB AB_5_65 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_65),
       .start_in   (start_in_5_65),
       .op_in      (op_in_5_65),
       .pivot_in   (pivot_in_5_65),
       .start_out  (start_out_5_65),
       .data_out   (data_out_5_65),
       .op_out     (op_out_5_65),
       .pivot_out  (pivot_out_5_65),
       .r          (r_5_65)
     );

  // row 5, col 66

     reg start_in_5_66;
     wire start_out_5_66;

     reg [1:0] op_in_5_66;
     wire [1:0] op_out_5_66;

     wire r_5_66;

     reg data_in_5_66;
     wire data_out_5_66;

     reg pivot_in_5_66;
     wire pivot_out_5_66;

     always @(posedge clk) begin
         op_in_5_66 <= op_out_5_65;
         pivot_in_5_66 <= pivot_out_5_65;
         start_in_5_66 <= start_out_5_65;
     end

     always @(posedge clk) begin
         data_in_5_66 <= data_out_4_66;
     end
  
     processor_AB AB_5_66 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_66),
       .start_in   (start_in_5_66),
       .op_in      (op_in_5_66),
       .pivot_in   (pivot_in_5_66),
       .start_out  (start_out_5_66),
       .data_out   (data_out_5_66),
       .op_out     (op_out_5_66),
       .pivot_out  (pivot_out_5_66),
       .r          (r_5_66)
     );

  // row 5, col 67

     reg start_in_5_67;
     wire start_out_5_67;

     reg [1:0] op_in_5_67;
     wire [1:0] op_out_5_67;

     wire r_5_67;

     reg data_in_5_67;
     wire data_out_5_67;

     reg pivot_in_5_67;
     wire pivot_out_5_67;

     always @(posedge clk) begin
         op_in_5_67 <= op_out_5_66;
         pivot_in_5_67 <= pivot_out_5_66;
         start_in_5_67 <= start_out_5_66;
     end

     always @(posedge clk) begin
         data_in_5_67 <= data_out_4_67;
     end
  
     processor_AB AB_5_67 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_67),
       .start_in   (start_in_5_67),
       .op_in      (op_in_5_67),
       .pivot_in   (pivot_in_5_67),
       .start_out  (start_out_5_67),
       .data_out   (data_out_5_67),
       .op_out     (op_out_5_67),
       .pivot_out  (pivot_out_5_67),
       .r          (r_5_67)
     );

  // row 5, col 68

     reg start_in_5_68;
     wire start_out_5_68;

     reg [1:0] op_in_5_68;
     wire [1:0] op_out_5_68;

     wire r_5_68;

     reg data_in_5_68;
     wire data_out_5_68;

     reg pivot_in_5_68;
     wire pivot_out_5_68;

     always @(posedge clk) begin
         op_in_5_68 <= op_out_5_67;
         pivot_in_5_68 <= pivot_out_5_67;
         start_in_5_68 <= start_out_5_67;
     end

     always @(posedge clk) begin
         data_in_5_68 <= data_out_4_68;
     end
  
     processor_AB AB_5_68 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_68),
       .start_in   (start_in_5_68),
       .op_in      (op_in_5_68),
       .pivot_in   (pivot_in_5_68),
       .start_out  (start_out_5_68),
       .data_out   (data_out_5_68),
       .op_out     (op_out_5_68),
       .pivot_out  (pivot_out_5_68),
       .r          (r_5_68)
     );

  // row 5, col 69

     reg start_in_5_69;
     wire start_out_5_69;

     reg [1:0] op_in_5_69;
     wire [1:0] op_out_5_69;

     wire r_5_69;

     reg data_in_5_69;
     wire data_out_5_69;

     reg pivot_in_5_69;
     wire pivot_out_5_69;

     always @(posedge clk) begin
         op_in_5_69 <= op_out_5_68;
         pivot_in_5_69 <= pivot_out_5_68;
         start_in_5_69 <= start_out_5_68;
     end

     always @(posedge clk) begin
         data_in_5_69 <= data_out_4_69;
     end
  
     processor_AB AB_5_69 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_69),
       .start_in   (start_in_5_69),
       .op_in      (op_in_5_69),
       .pivot_in   (pivot_in_5_69),
       .start_out  (start_out_5_69),
       .data_out   (data_out_5_69),
       .op_out     (op_out_5_69),
       .pivot_out  (pivot_out_5_69),
       .r          (r_5_69)
     );

  // row 5, col 70

     reg start_in_5_70;
     wire start_out_5_70;

     reg [1:0] op_in_5_70;
     wire [1:0] op_out_5_70;

     wire r_5_70;

     reg data_in_5_70;
     wire data_out_5_70;

     reg pivot_in_5_70;
     wire pivot_out_5_70;

     always @(posedge clk) begin
         op_in_5_70 <= op_out_5_69;
         pivot_in_5_70 <= pivot_out_5_69;
         start_in_5_70 <= start_out_5_69;
     end

     always @(posedge clk) begin
         data_in_5_70 <= data_out_4_70;
     end
  
     processor_AB AB_5_70 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_70),
       .start_in   (start_in_5_70),
       .op_in      (op_in_5_70),
       .pivot_in   (pivot_in_5_70),
       .start_out  (start_out_5_70),
       .data_out   (data_out_5_70),
       .op_out     (op_out_5_70),
       .pivot_out  (pivot_out_5_70),
       .r          (r_5_70)
     );

  // row 5, col 71

     reg start_in_5_71;
     wire start_out_5_71;

     reg [1:0] op_in_5_71;
     wire [1:0] op_out_5_71;

     wire r_5_71;

     reg data_in_5_71;
     wire data_out_5_71;

     reg pivot_in_5_71;
     wire pivot_out_5_71;

     always @(posedge clk) begin
         op_in_5_71 <= op_out_5_70;
         pivot_in_5_71 <= pivot_out_5_70;
         start_in_5_71 <= start_out_5_70;
     end

     always @(posedge clk) begin
         data_in_5_71 <= data_out_4_71;
     end
  
     processor_AB AB_5_71 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_71),
       .start_in   (start_in_5_71),
       .op_in      (op_in_5_71),
       .pivot_in   (pivot_in_5_71),
       .start_out  (start_out_5_71),
       .data_out   (data_out_5_71),
       .op_out     (op_out_5_71),
       .pivot_out  (pivot_out_5_71),
       .r          (r_5_71)
     );

  // row 5, col 72

     reg start_in_5_72;
     wire start_out_5_72;

     reg [1:0] op_in_5_72;
     wire [1:0] op_out_5_72;

     wire r_5_72;

     reg data_in_5_72;
     wire data_out_5_72;

     reg pivot_in_5_72;
     wire pivot_out_5_72;

     always @(posedge clk) begin
         op_in_5_72 <= op_out_5_71;
         pivot_in_5_72 <= pivot_out_5_71;
         start_in_5_72 <= start_out_5_71;
     end

     always @(posedge clk) begin
         data_in_5_72 <= data_out_4_72;
     end
  
     processor_AB AB_5_72 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_72),
       .start_in   (start_in_5_72),
       .op_in      (op_in_5_72),
       .pivot_in   (pivot_in_5_72),
       .start_out  (start_out_5_72),
       .data_out   (data_out_5_72),
       .op_out     (op_out_5_72),
       .pivot_out  (pivot_out_5_72),
       .r          (r_5_72)
     );

  // row 5, col 73

     reg start_in_5_73;
     wire start_out_5_73;

     reg [1:0] op_in_5_73;
     wire [1:0] op_out_5_73;

     wire r_5_73;

     reg data_in_5_73;
     wire data_out_5_73;

     reg pivot_in_5_73;
     wire pivot_out_5_73;

     always @(posedge clk) begin
         op_in_5_73 <= op_out_5_72;
         pivot_in_5_73 <= pivot_out_5_72;
         start_in_5_73 <= start_out_5_72;
     end

     always @(posedge clk) begin
         data_in_5_73 <= data_out_4_73;
     end
  
     processor_AB AB_5_73 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_73),
       .start_in   (start_in_5_73),
       .op_in      (op_in_5_73),
       .pivot_in   (pivot_in_5_73),
       .start_out  (start_out_5_73),
       .data_out   (data_out_5_73),
       .op_out     (op_out_5_73),
       .pivot_out  (pivot_out_5_73),
       .r          (r_5_73)
     );

  // row 5, col 74

     reg start_in_5_74;
     wire start_out_5_74;

     reg [1:0] op_in_5_74;
     wire [1:0] op_out_5_74;

     wire r_5_74;

     reg data_in_5_74;
     wire data_out_5_74;

     reg pivot_in_5_74;
     wire pivot_out_5_74;

     always @(posedge clk) begin
         op_in_5_74 <= op_out_5_73;
         pivot_in_5_74 <= pivot_out_5_73;
         start_in_5_74 <= start_out_5_73;
     end

     always @(posedge clk) begin
         data_in_5_74 <= data_out_4_74;
     end
  
     processor_AB AB_5_74 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_74),
       .start_in   (start_in_5_74),
       .op_in      (op_in_5_74),
       .pivot_in   (pivot_in_5_74),
       .start_out  (start_out_5_74),
       .data_out   (data_out_5_74),
       .op_out     (op_out_5_74),
       .pivot_out  (pivot_out_5_74),
       .r          (r_5_74)
     );

  // row 5, col 75

     reg start_in_5_75;
     wire start_out_5_75;

     reg [1:0] op_in_5_75;
     wire [1:0] op_out_5_75;

     wire r_5_75;

     reg data_in_5_75;
     wire data_out_5_75;

     reg pivot_in_5_75;
     wire pivot_out_5_75;

     always @(posedge clk) begin
         op_in_5_75 <= op_out_5_74;
         pivot_in_5_75 <= pivot_out_5_74;
         start_in_5_75 <= start_out_5_74;
     end

     always @(posedge clk) begin
         data_in_5_75 <= data_out_4_75;
     end
  
     processor_AB AB_5_75 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_75),
       .start_in   (start_in_5_75),
       .op_in      (op_in_5_75),
       .pivot_in   (pivot_in_5_75),
       .start_out  (start_out_5_75),
       .data_out   (data_out_5_75),
       .op_out     (op_out_5_75),
       .pivot_out  (pivot_out_5_75),
       .r          (r_5_75)
     );

  // row 5, col 76

     reg start_in_5_76;
     wire start_out_5_76;

     reg [1:0] op_in_5_76;
     wire [1:0] op_out_5_76;

     wire r_5_76;

     reg data_in_5_76;
     wire data_out_5_76;

     reg pivot_in_5_76;
     wire pivot_out_5_76;

     always @(posedge clk) begin
         op_in_5_76 <= op_out_5_75;
         pivot_in_5_76 <= pivot_out_5_75;
         start_in_5_76 <= start_out_5_75;
     end

     always @(posedge clk) begin
         data_in_5_76 <= data_out_4_76;
     end
  
     processor_AB AB_5_76 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_76),
       .start_in   (start_in_5_76),
       .op_in      (op_in_5_76),
       .pivot_in   (pivot_in_5_76),
       .start_out  (start_out_5_76),
       .data_out   (data_out_5_76),
       .op_out     (op_out_5_76),
       .pivot_out  (pivot_out_5_76),
       .r          (r_5_76)
     );

  // row 5, col 77

     reg start_in_5_77;
     wire start_out_5_77;

     reg [1:0] op_in_5_77;
     wire [1:0] op_out_5_77;

     wire r_5_77;

     reg data_in_5_77;
     wire data_out_5_77;

     reg pivot_in_5_77;
     wire pivot_out_5_77;

     always @(posedge clk) begin
         op_in_5_77 <= op_out_5_76;
         pivot_in_5_77 <= pivot_out_5_76;
         start_in_5_77 <= start_out_5_76;
     end

     always @(posedge clk) begin
         data_in_5_77 <= data_out_4_77;
     end
  
     processor_AB AB_5_77 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_77),
       .start_in   (start_in_5_77),
       .op_in      (op_in_5_77),
       .pivot_in   (pivot_in_5_77),
       .start_out  (start_out_5_77),
       .data_out   (data_out_5_77),
       .op_out     (op_out_5_77),
       .pivot_out  (pivot_out_5_77),
       .r          (r_5_77)
     );

  // row 5, col 78

     reg start_in_5_78;
     wire start_out_5_78;

     reg [1:0] op_in_5_78;
     wire [1:0] op_out_5_78;

     wire r_5_78;

     reg data_in_5_78;
     wire data_out_5_78;

     reg pivot_in_5_78;
     wire pivot_out_5_78;

     always @(posedge clk) begin
         op_in_5_78 <= op_out_5_77;
         pivot_in_5_78 <= pivot_out_5_77;
         start_in_5_78 <= start_out_5_77;
     end

     always @(posedge clk) begin
         data_in_5_78 <= data_out_4_78;
     end
  
     processor_AB AB_5_78 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_78),
       .start_in   (start_in_5_78),
       .op_in      (op_in_5_78),
       .pivot_in   (pivot_in_5_78),
       .start_out  (start_out_5_78),
       .data_out   (data_out_5_78),
       .op_out     (op_out_5_78),
       .pivot_out  (pivot_out_5_78),
       .r          (r_5_78)
     );

  // row 5, col 79

     reg start_in_5_79;
     wire start_out_5_79;

     reg [1:0] op_in_5_79;
     wire [1:0] op_out_5_79;

     wire r_5_79;

     reg data_in_5_79;
     wire data_out_5_79;

     reg pivot_in_5_79;
     wire pivot_out_5_79;

     always @(posedge clk) begin
         op_in_5_79 <= op_out_5_78;
         pivot_in_5_79 <= pivot_out_5_78;
         start_in_5_79 <= start_out_5_78;
     end

     always @(posedge clk) begin
         data_in_5_79 <= data_out_4_79;
     end
  
     processor_AB AB_5_79 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_79),
       .start_in   (start_in_5_79),
       .op_in      (op_in_5_79),
       .pivot_in   (pivot_in_5_79),
       .start_out  (start_out_5_79),
       .data_out   (data_out_5_79),
       .op_out     (op_out_5_79),
       .pivot_out  (pivot_out_5_79),
       .r          (r_5_79)
     );

  // row 5, col 80

     reg start_in_5_80;
     wire start_out_5_80;

     reg [1:0] op_in_5_80;
     wire [1:0] op_out_5_80;

     wire r_5_80;

     reg data_in_5_80;
     wire data_out_5_80;

     reg pivot_in_5_80;
     wire pivot_out_5_80;

     always @(posedge clk) begin
         op_in_5_80 <= op_out_5_79;
         pivot_in_5_80 <= pivot_out_5_79;
         start_in_5_80 <= start_out_5_79;
     end

     always @(posedge clk) begin
         data_in_5_80 <= data_out_4_80;
     end
  
     processor_AB AB_5_80 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_80),
       .start_in   (start_in_5_80),
       .op_in      (op_in_5_80),
       .pivot_in   (pivot_in_5_80),
       .start_out  (start_out_5_80),
       .data_out   (data_out_5_80),
       .op_out     (op_out_5_80),
       .pivot_out  (pivot_out_5_80),
       .r          (r_5_80)
     );

  // row 5, col 81

     reg start_in_5_81;
     wire start_out_5_81;

     reg [1:0] op_in_5_81;
     wire [1:0] op_out_5_81;

     wire r_5_81;

     reg data_in_5_81;
     wire data_out_5_81;

     reg pivot_in_5_81;
     wire pivot_out_5_81;

     always @(posedge clk) begin
         op_in_5_81 <= op_out_5_80;
         pivot_in_5_81 <= pivot_out_5_80;
         start_in_5_81 <= start_out_5_80;
     end

     always @(posedge clk) begin
         data_in_5_81 <= data_out_4_81;
     end
  
     processor_AB AB_5_81 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_81),
       .start_in   (start_in_5_81),
       .op_in      (op_in_5_81),
       .pivot_in   (pivot_in_5_81),
       .start_out  (start_out_5_81),
       .data_out   (data_out_5_81),
       .op_out     (op_out_5_81),
       .pivot_out  (pivot_out_5_81),
       .r          (r_5_81)
     );

  // row 5, col 82

     reg start_in_5_82;
     wire start_out_5_82;

     reg [1:0] op_in_5_82;
     wire [1:0] op_out_5_82;

     wire r_5_82;

     reg data_in_5_82;
     wire data_out_5_82;

     reg pivot_in_5_82;
     wire pivot_out_5_82;

     always @(posedge clk) begin
         op_in_5_82 <= op_out_5_81;
         pivot_in_5_82 <= pivot_out_5_81;
         start_in_5_82 <= start_out_5_81;
     end

     always @(posedge clk) begin
         data_in_5_82 <= data_out_4_82;
     end
  
     processor_AB AB_5_82 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_82),
       .start_in   (start_in_5_82),
       .op_in      (op_in_5_82),
       .pivot_in   (pivot_in_5_82),
       .start_out  (start_out_5_82),
       .data_out   (data_out_5_82),
       .op_out     (op_out_5_82),
       .pivot_out  (pivot_out_5_82),
       .r          (r_5_82)
     );

  // row 5, col 83

     reg start_in_5_83;
     wire start_out_5_83;

     reg [1:0] op_in_5_83;
     wire [1:0] op_out_5_83;

     wire r_5_83;

     reg data_in_5_83;
     wire data_out_5_83;

     reg pivot_in_5_83;
     wire pivot_out_5_83;

     always @(posedge clk) begin
         op_in_5_83 <= op_out_5_82;
         pivot_in_5_83 <= pivot_out_5_82;
         start_in_5_83 <= start_out_5_82;
     end

     always @(posedge clk) begin
         data_in_5_83 <= data_out_4_83;
     end
  
     processor_AB AB_5_83 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_83),
       .start_in   (start_in_5_83),
       .op_in      (op_in_5_83),
       .pivot_in   (pivot_in_5_83),
       .start_out  (start_out_5_83),
       .data_out   (data_out_5_83),
       .op_out     (op_out_5_83),
       .pivot_out  (pivot_out_5_83),
       .r          (r_5_83)
     );

  // row 5, col 84

     reg start_in_5_84;
     wire start_out_5_84;

     reg [1:0] op_in_5_84;
     wire [1:0] op_out_5_84;

     wire r_5_84;

     reg data_in_5_84;
     wire data_out_5_84;

     reg pivot_in_5_84;
     wire pivot_out_5_84;

     always @(posedge clk) begin
         op_in_5_84 <= op_out_5_83;
         pivot_in_5_84 <= pivot_out_5_83;
         start_in_5_84 <= start_out_5_83;
     end

     always @(posedge clk) begin
         data_in_5_84 <= data_out_4_84;
     end
  
     processor_AB AB_5_84 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_84),
       .start_in   (start_in_5_84),
       .op_in      (op_in_5_84),
       .pivot_in   (pivot_in_5_84),
       .start_out  (start_out_5_84),
       .data_out   (data_out_5_84),
       .op_out     (op_out_5_84),
       .pivot_out  (pivot_out_5_84),
       .r          (r_5_84)
     );

  // row 5, col 85

     reg start_in_5_85;
     wire start_out_5_85;

     reg [1:0] op_in_5_85;
     wire [1:0] op_out_5_85;

     wire r_5_85;

     reg data_in_5_85;
     wire data_out_5_85;

     reg pivot_in_5_85;
     wire pivot_out_5_85;

     always @(posedge clk) begin
         op_in_5_85 <= op_out_5_84;
         pivot_in_5_85 <= pivot_out_5_84;
         start_in_5_85 <= start_out_5_84;
     end

     always @(posedge clk) begin
         data_in_5_85 <= data_out_4_85;
     end
  
     processor_AB AB_5_85 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_85),
       .start_in   (start_in_5_85),
       .op_in      (op_in_5_85),
       .pivot_in   (pivot_in_5_85),
       .start_out  (start_out_5_85),
       .data_out   (data_out_5_85),
       .op_out     (op_out_5_85),
       .pivot_out  (pivot_out_5_85),
       .r          (r_5_85)
     );

  // row 5, col 86

     reg start_in_5_86;
     wire start_out_5_86;

     reg [1:0] op_in_5_86;
     wire [1:0] op_out_5_86;

     wire r_5_86;

     reg data_in_5_86;
     wire data_out_5_86;

     reg pivot_in_5_86;
     wire pivot_out_5_86;

     always @(posedge clk) begin
         op_in_5_86 <= op_out_5_85;
         pivot_in_5_86 <= pivot_out_5_85;
         start_in_5_86 <= start_out_5_85;
     end

     always @(posedge clk) begin
         data_in_5_86 <= data_out_4_86;
     end
  
     processor_AB AB_5_86 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_86),
       .start_in   (start_in_5_86),
       .op_in      (op_in_5_86),
       .pivot_in   (pivot_in_5_86),
       .start_out  (start_out_5_86),
       .data_out   (data_out_5_86),
       .op_out     (op_out_5_86),
       .pivot_out  (pivot_out_5_86),
       .r          (r_5_86)
     );

  // row 5, col 87

     reg start_in_5_87;
     wire start_out_5_87;

     reg [1:0] op_in_5_87;
     wire [1:0] op_out_5_87;

     wire r_5_87;

     reg data_in_5_87;
     wire data_out_5_87;

     reg pivot_in_5_87;
     wire pivot_out_5_87;

     always @(posedge clk) begin
         op_in_5_87 <= op_out_5_86;
         pivot_in_5_87 <= pivot_out_5_86;
         start_in_5_87 <= start_out_5_86;
     end

     always @(posedge clk) begin
         data_in_5_87 <= data_out_4_87;
     end
  
     processor_AB AB_5_87 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_87),
       .start_in   (start_in_5_87),
       .op_in      (op_in_5_87),
       .pivot_in   (pivot_in_5_87),
       .start_out  (start_out_5_87),
       .data_out   (data_out_5_87),
       .op_out     (op_out_5_87),
       .pivot_out  (pivot_out_5_87),
       .r          (r_5_87)
     );

  // row 5, col 88

     reg start_in_5_88;
     wire start_out_5_88;

     reg [1:0] op_in_5_88;
     wire [1:0] op_out_5_88;

     wire r_5_88;

     reg data_in_5_88;
     wire data_out_5_88;

     reg pivot_in_5_88;
     wire pivot_out_5_88;

     always @(posedge clk) begin
         op_in_5_88 <= op_out_5_87;
         pivot_in_5_88 <= pivot_out_5_87;
         start_in_5_88 <= start_out_5_87;
     end

     always @(posedge clk) begin
         data_in_5_88 <= data_out_4_88;
     end
  
     processor_AB AB_5_88 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_88),
       .start_in   (start_in_5_88),
       .op_in      (op_in_5_88),
       .pivot_in   (pivot_in_5_88),
       .start_out  (start_out_5_88),
       .data_out   (data_out_5_88),
       .op_out     (op_out_5_88),
       .pivot_out  (pivot_out_5_88),
       .r          (r_5_88)
     );

  // row 5, col 89

     reg start_in_5_89;
     wire start_out_5_89;

     reg [1:0] op_in_5_89;
     wire [1:0] op_out_5_89;

     wire r_5_89;

     reg data_in_5_89;
     wire data_out_5_89;

     reg pivot_in_5_89;
     wire pivot_out_5_89;

     always @(posedge clk) begin
         op_in_5_89 <= op_out_5_88;
         pivot_in_5_89 <= pivot_out_5_88;
         start_in_5_89 <= start_out_5_88;
     end

     always @(posedge clk) begin
         data_in_5_89 <= data_out_4_89;
     end
  
     processor_AB AB_5_89 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_89),
       .start_in   (start_in_5_89),
       .op_in      (op_in_5_89),
       .pivot_in   (pivot_in_5_89),
       .start_out  (start_out_5_89),
       .data_out   (data_out_5_89),
       .op_out     (op_out_5_89),
       .pivot_out  (pivot_out_5_89),
       .r          (r_5_89)
     );

  // row 5, col 90

     reg start_in_5_90;
     wire start_out_5_90;

     reg [1:0] op_in_5_90;
     wire [1:0] op_out_5_90;

     wire r_5_90;

     reg data_in_5_90;
     wire data_out_5_90;

     reg pivot_in_5_90;
     wire pivot_out_5_90;

     always @(posedge clk) begin
         op_in_5_90 <= op_out_5_89;
         pivot_in_5_90 <= pivot_out_5_89;
         start_in_5_90 <= start_out_5_89;
     end

     always @(posedge clk) begin
         data_in_5_90 <= data_out_4_90;
     end
  
     processor_AB AB_5_90 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_90),
       .start_in   (start_in_5_90),
       .op_in      (op_in_5_90),
       .pivot_in   (pivot_in_5_90),
       .start_out  (start_out_5_90),
       .data_out   (data_out_5_90),
       .op_out     (op_out_5_90),
       .pivot_out  (pivot_out_5_90),
       .r          (r_5_90)
     );

  // row 5, col 91

     reg start_in_5_91;
     wire start_out_5_91;

     reg [1:0] op_in_5_91;
     wire [1:0] op_out_5_91;

     wire r_5_91;

     reg data_in_5_91;
     wire data_out_5_91;

     reg pivot_in_5_91;
     wire pivot_out_5_91;

     always @(posedge clk) begin
         op_in_5_91 <= op_out_5_90;
         pivot_in_5_91 <= pivot_out_5_90;
         start_in_5_91 <= start_out_5_90;
     end

     always @(posedge clk) begin
         data_in_5_91 <= data_out_4_91;
     end
  
     processor_AB AB_5_91 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_91),
       .start_in   (start_in_5_91),
       .op_in      (op_in_5_91),
       .pivot_in   (pivot_in_5_91),
       .start_out  (start_out_5_91),
       .data_out   (data_out_5_91),
       .op_out     (op_out_5_91),
       .pivot_out  (pivot_out_5_91),
       .r          (r_5_91)
     );

  // row 5, col 92

     reg start_in_5_92;
     wire start_out_5_92;

     reg [1:0] op_in_5_92;
     wire [1:0] op_out_5_92;

     wire r_5_92;

     reg data_in_5_92;
     wire data_out_5_92;

     reg pivot_in_5_92;
     wire pivot_out_5_92;

     always @(posedge clk) begin
         op_in_5_92 <= op_out_5_91;
         pivot_in_5_92 <= pivot_out_5_91;
         start_in_5_92 <= start_out_5_91;
     end

     always @(posedge clk) begin
         data_in_5_92 <= data_out_4_92;
     end
  
     processor_AB AB_5_92 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_92),
       .start_in   (start_in_5_92),
       .op_in      (op_in_5_92),
       .pivot_in   (pivot_in_5_92),
       .start_out  (start_out_5_92),
       .data_out   (data_out_5_92),
       .op_out     (op_out_5_92),
       .pivot_out  (pivot_out_5_92),
       .r          (r_5_92)
     );

  // row 5, col 93

     reg start_in_5_93;
     wire start_out_5_93;

     reg [1:0] op_in_5_93;
     wire [1:0] op_out_5_93;

     wire r_5_93;

     reg data_in_5_93;
     wire data_out_5_93;

     reg pivot_in_5_93;
     wire pivot_out_5_93;

     always @(posedge clk) begin
         op_in_5_93 <= op_out_5_92;
         pivot_in_5_93 <= pivot_out_5_92;
         start_in_5_93 <= start_out_5_92;
     end

     always @(posedge clk) begin
         data_in_5_93 <= data_out_4_93;
     end
  
     processor_AB AB_5_93 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_93),
       .start_in   (start_in_5_93),
       .op_in      (op_in_5_93),
       .pivot_in   (pivot_in_5_93),
       .start_out  (start_out_5_93),
       .data_out   (data_out_5_93),
       .op_out     (op_out_5_93),
       .pivot_out  (pivot_out_5_93),
       .r          (r_5_93)
     );

  // row 5, col 94

     reg start_in_5_94;
     wire start_out_5_94;

     reg [1:0] op_in_5_94;
     wire [1:0] op_out_5_94;

     wire r_5_94;

     reg data_in_5_94;
     wire data_out_5_94;

     reg pivot_in_5_94;
     wire pivot_out_5_94;

     always @(posedge clk) begin
         op_in_5_94 <= op_out_5_93;
         pivot_in_5_94 <= pivot_out_5_93;
         start_in_5_94 <= start_out_5_93;
     end

     always @(posedge clk) begin
         data_in_5_94 <= data_out_4_94;
     end
  
     processor_AB AB_5_94 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_94),
       .start_in   (start_in_5_94),
       .op_in      (op_in_5_94),
       .pivot_in   (pivot_in_5_94),
       .start_out  (start_out_5_94),
       .data_out   (data_out_5_94),
       .op_out     (op_out_5_94),
       .pivot_out  (pivot_out_5_94),
       .r          (r_5_94)
     );

  // row 5, col 95

     reg start_in_5_95;
     wire start_out_5_95;

     reg [1:0] op_in_5_95;
     wire [1:0] op_out_5_95;

     wire r_5_95;

     reg data_in_5_95;
     wire data_out_5_95;

     reg pivot_in_5_95;
     wire pivot_out_5_95;

     always @(posedge clk) begin
         op_in_5_95 <= op_out_5_94;
         pivot_in_5_95 <= pivot_out_5_94;
         start_in_5_95 <= start_out_5_94;
     end

     always @(posedge clk) begin
         data_in_5_95 <= data_out_4_95;
     end
  
     processor_AB AB_5_95 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_95),
       .start_in   (start_in_5_95),
       .op_in      (op_in_5_95),
       .pivot_in   (pivot_in_5_95),
       .start_out  (start_out_5_95),
       .data_out   (data_out_5_95),
       .op_out     (op_out_5_95),
       .pivot_out  (pivot_out_5_95),
       .r          (r_5_95)
     );

  // row 5, col 96

     reg start_in_5_96;
     wire start_out_5_96;

     reg [1:0] op_in_5_96;
     wire [1:0] op_out_5_96;

     wire r_5_96;

     reg data_in_5_96;
     wire data_out_5_96;

     reg pivot_in_5_96;
     wire pivot_out_5_96;

     always @(posedge clk) begin
         op_in_5_96 <= op_out_5_95;
         pivot_in_5_96 <= pivot_out_5_95;
         start_in_5_96 <= start_out_5_95;
     end

     always @(posedge clk) begin
         data_in_5_96 <= data_out_4_96;
     end
  
     processor_AB AB_5_96 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_96),
       .start_in   (start_in_5_96),
       .op_in      (op_in_5_96),
       .pivot_in   (pivot_in_5_96),
       .start_out  (start_out_5_96),
       .data_out   (data_out_5_96),
       .op_out     (op_out_5_96),
       .pivot_out  (pivot_out_5_96),
       .r          (r_5_96)
     );

  // row 5, col 97

     reg start_in_5_97;
     wire start_out_5_97;

     reg [1:0] op_in_5_97;
     wire [1:0] op_out_5_97;

     wire r_5_97;

     reg data_in_5_97;
     wire data_out_5_97;

     reg pivot_in_5_97;
     wire pivot_out_5_97;

     always @(posedge clk) begin
         op_in_5_97 <= op_out_5_96;
         pivot_in_5_97 <= pivot_out_5_96;
         start_in_5_97 <= start_out_5_96;
     end

     always @(posedge clk) begin
         data_in_5_97 <= data_out_4_97;
     end
  
     processor_AB AB_5_97 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_97),
       .start_in   (start_in_5_97),
       .op_in      (op_in_5_97),
       .pivot_in   (pivot_in_5_97),
       .start_out  (start_out_5_97),
       .data_out   (data_out_5_97),
       .op_out     (op_out_5_97),
       .pivot_out  (pivot_out_5_97),
       .r          (r_5_97)
     );

  // row 5, col 98

     reg start_in_5_98;
     wire start_out_5_98;

     reg [1:0] op_in_5_98;
     wire [1:0] op_out_5_98;

     wire r_5_98;

     reg data_in_5_98;
     wire data_out_5_98;

     reg pivot_in_5_98;
     wire pivot_out_5_98;

     always @(posedge clk) begin
         op_in_5_98 <= op_out_5_97;
         pivot_in_5_98 <= pivot_out_5_97;
         start_in_5_98 <= start_out_5_97;
     end

     always @(posedge clk) begin
         data_in_5_98 <= data_out_4_98;
     end
  
     processor_AB AB_5_98 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_98),
       .start_in   (start_in_5_98),
       .op_in      (op_in_5_98),
       .pivot_in   (pivot_in_5_98),
       .start_out  (start_out_5_98),
       .data_out   (data_out_5_98),
       .op_out     (op_out_5_98),
       .pivot_out  (pivot_out_5_98),
       .r          (r_5_98)
     );

  // row 5, col 99

     reg start_in_5_99;
     wire start_out_5_99;

     reg [1:0] op_in_5_99;
     wire [1:0] op_out_5_99;

     wire r_5_99;

     reg data_in_5_99;
     wire data_out_5_99;

     reg pivot_in_5_99;
     wire pivot_out_5_99;

     always @(posedge clk) begin
         op_in_5_99 <= op_out_5_98;
         pivot_in_5_99 <= pivot_out_5_98;
         start_in_5_99 <= start_out_5_98;
     end

     always @(posedge clk) begin
         data_in_5_99 <= data_out_4_99;
     end
  
     processor_AB AB_5_99 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_99),
       .start_in   (start_in_5_99),
       .op_in      (op_in_5_99),
       .pivot_in   (pivot_in_5_99),
       .start_out  (start_out_5_99),
       .data_out   (data_out_5_99),
       .op_out     (op_out_5_99),
       .pivot_out  (pivot_out_5_99),
       .r          (r_5_99)
     );

  // row 5, col 100

     reg start_in_5_100;
     wire start_out_5_100;

     reg [1:0] op_in_5_100;
     wire [1:0] op_out_5_100;

     wire r_5_100;

     reg data_in_5_100;
     wire data_out_5_100;

     reg pivot_in_5_100;
     wire pivot_out_5_100;

     always @(posedge clk) begin
         op_in_5_100 <= op_out_5_99;
         pivot_in_5_100 <= pivot_out_5_99;
         start_in_5_100 <= start_out_5_99;
     end

     always @(posedge clk) begin
         data_in_5_100 <= data_out_4_100;
     end
  
     processor_AB AB_5_100 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_5_100),
       .start_in   (start_in_5_100),
       .op_in      (op_in_5_100),
       .pivot_in   (pivot_in_5_100),
       .start_out  (start_out_5_100),
       .data_out   (data_out_5_100),
       .op_out     (op_out_5_100),
       .pivot_out  (pivot_out_5_100),
       .r          (r_5_100)
     );

  /////////////////////////////////////
  // outputs 

  wire [5:0] pivot_found;
  wire [100:0] row0, row1, row2, row3, row4, row5;

  assign pivot_found = {r_0_0 | r_0_1 | r_0_2 | r_0_3 | r_0_4 | r_0_5 | r_0_6 | r_0_7 | r_0_8 | r_0_9 | r_0_10 | r_0_11 | r_0_12 | r_0_13 | r_0_14 | r_0_15 | r_0_16 | r_0_17 | r_0_18 | r_0_19 | r_0_20 | r_0_21 | r_0_22 | r_0_23 | r_0_24 | r_0_25 | r_0_26 | r_0_27 | r_0_28 | r_0_29 | r_0_30 | r_0_31 | r_0_32 | r_0_33 | r_0_34 | r_0_35 | r_0_36 | r_0_37 | r_0_38 | r_0_39 | r_0_40 | r_0_41 | r_0_42 | r_0_43 | r_0_44 | r_0_45 | r_0_46 | r_0_47 | r_0_48 | r_0_49 | r_0_50 | r_0_51 | r_0_52 | r_0_53 | r_0_54 | r_0_55 | r_0_56 | r_0_57 | r_0_58 | r_0_59 | r_0_60 | r_0_61 | r_0_62 | r_0_63 | r_0_64 | r_0_65 | r_0_66 | r_0_67 | r_0_68 | r_0_69 | r_0_70 | r_0_71 | r_0_72 | r_0_73 | r_0_74 | r_0_75 | r_0_76 | r_0_77 | r_0_78 | r_0_79 | r_0_80 | r_0_81 | r_0_82 | r_0_83 | r_0_84 | r_0_85 | r_0_86 | r_0_87 | r_0_88 | r_0_89 | r_0_90 | r_0_91 | r_0_92 | r_0_93 | r_0_94 | r_0_95 | r_0_96 | r_0_97 | r_0_98 | r_0_99 | r_0_100, r_1_0 | r_1_1 | r_1_2 | r_1_3 | r_1_4 | r_1_5 | r_1_6 | r_1_7 | r_1_8 | r_1_9 | r_1_10 | r_1_11 | r_1_12 | r_1_13 | r_1_14 | r_1_15 | r_1_16 | r_1_17 | r_1_18 | r_1_19 | r_1_20 | r_1_21 | r_1_22 | r_1_23 | r_1_24 | r_1_25 | r_1_26 | r_1_27 | r_1_28 | r_1_29 | r_1_30 | r_1_31 | r_1_32 | r_1_33 | r_1_34 | r_1_35 | r_1_36 | r_1_37 | r_1_38 | r_1_39 | r_1_40 | r_1_41 | r_1_42 | r_1_43 | r_1_44 | r_1_45 | r_1_46 | r_1_47 | r_1_48 | r_1_49 | r_1_50 | r_1_51 | r_1_52 | r_1_53 | r_1_54 | r_1_55 | r_1_56 | r_1_57 | r_1_58 | r_1_59 | r_1_60 | r_1_61 | r_1_62 | r_1_63 | r_1_64 | r_1_65 | r_1_66 | r_1_67 | r_1_68 | r_1_69 | r_1_70 | r_1_71 | r_1_72 | r_1_73 | r_1_74 | r_1_75 | r_1_76 | r_1_77 | r_1_78 | r_1_79 | r_1_80 | r_1_81 | r_1_82 | r_1_83 | r_1_84 | r_1_85 | r_1_86 | r_1_87 | r_1_88 | r_1_89 | r_1_90 | r_1_91 | r_1_92 | r_1_93 | r_1_94 | r_1_95 | r_1_96 | r_1_97 | r_1_98 | r_1_99 | r_1_100, r_2_0 | r_2_1 | r_2_2 | r_2_3 | r_2_4 | r_2_5 | r_2_6 | r_2_7 | r_2_8 | r_2_9 | r_2_10 | r_2_11 | r_2_12 | r_2_13 | r_2_14 | r_2_15 | r_2_16 | r_2_17 | r_2_18 | r_2_19 | r_2_20 | r_2_21 | r_2_22 | r_2_23 | r_2_24 | r_2_25 | r_2_26 | r_2_27 | r_2_28 | r_2_29 | r_2_30 | r_2_31 | r_2_32 | r_2_33 | r_2_34 | r_2_35 | r_2_36 | r_2_37 | r_2_38 | r_2_39 | r_2_40 | r_2_41 | r_2_42 | r_2_43 | r_2_44 | r_2_45 | r_2_46 | r_2_47 | r_2_48 | r_2_49 | r_2_50 | r_2_51 | r_2_52 | r_2_53 | r_2_54 | r_2_55 | r_2_56 | r_2_57 | r_2_58 | r_2_59 | r_2_60 | r_2_61 | r_2_62 | r_2_63 | r_2_64 | r_2_65 | r_2_66 | r_2_67 | r_2_68 | r_2_69 | r_2_70 | r_2_71 | r_2_72 | r_2_73 | r_2_74 | r_2_75 | r_2_76 | r_2_77 | r_2_78 | r_2_79 | r_2_80 | r_2_81 | r_2_82 | r_2_83 | r_2_84 | r_2_85 | r_2_86 | r_2_87 | r_2_88 | r_2_89 | r_2_90 | r_2_91 | r_2_92 | r_2_93 | r_2_94 | r_2_95 | r_2_96 | r_2_97 | r_2_98 | r_2_99 | r_2_100, r_3_0 | r_3_1 | r_3_2 | r_3_3 | r_3_4 | r_3_5 | r_3_6 | r_3_7 | r_3_8 | r_3_9 | r_3_10 | r_3_11 | r_3_12 | r_3_13 | r_3_14 | r_3_15 | r_3_16 | r_3_17 | r_3_18 | r_3_19 | r_3_20 | r_3_21 | r_3_22 | r_3_23 | r_3_24 | r_3_25 | r_3_26 | r_3_27 | r_3_28 | r_3_29 | r_3_30 | r_3_31 | r_3_32 | r_3_33 | r_3_34 | r_3_35 | r_3_36 | r_3_37 | r_3_38 | r_3_39 | r_3_40 | r_3_41 | r_3_42 | r_3_43 | r_3_44 | r_3_45 | r_3_46 | r_3_47 | r_3_48 | r_3_49 | r_3_50 | r_3_51 | r_3_52 | r_3_53 | r_3_54 | r_3_55 | r_3_56 | r_3_57 | r_3_58 | r_3_59 | r_3_60 | r_3_61 | r_3_62 | r_3_63 | r_3_64 | r_3_65 | r_3_66 | r_3_67 | r_3_68 | r_3_69 | r_3_70 | r_3_71 | r_3_72 | r_3_73 | r_3_74 | r_3_75 | r_3_76 | r_3_77 | r_3_78 | r_3_79 | r_3_80 | r_3_81 | r_3_82 | r_3_83 | r_3_84 | r_3_85 | r_3_86 | r_3_87 | r_3_88 | r_3_89 | r_3_90 | r_3_91 | r_3_92 | r_3_93 | r_3_94 | r_3_95 | r_3_96 | r_3_97 | r_3_98 | r_3_99 | r_3_100, r_4_0 | r_4_1 | r_4_2 | r_4_3 | r_4_4 | r_4_5 | r_4_6 | r_4_7 | r_4_8 | r_4_9 | r_4_10 | r_4_11 | r_4_12 | r_4_13 | r_4_14 | r_4_15 | r_4_16 | r_4_17 | r_4_18 | r_4_19 | r_4_20 | r_4_21 | r_4_22 | r_4_23 | r_4_24 | r_4_25 | r_4_26 | r_4_27 | r_4_28 | r_4_29 | r_4_30 | r_4_31 | r_4_32 | r_4_33 | r_4_34 | r_4_35 | r_4_36 | r_4_37 | r_4_38 | r_4_39 | r_4_40 | r_4_41 | r_4_42 | r_4_43 | r_4_44 | r_4_45 | r_4_46 | r_4_47 | r_4_48 | r_4_49 | r_4_50 | r_4_51 | r_4_52 | r_4_53 | r_4_54 | r_4_55 | r_4_56 | r_4_57 | r_4_58 | r_4_59 | r_4_60 | r_4_61 | r_4_62 | r_4_63 | r_4_64 | r_4_65 | r_4_66 | r_4_67 | r_4_68 | r_4_69 | r_4_70 | r_4_71 | r_4_72 | r_4_73 | r_4_74 | r_4_75 | r_4_76 | r_4_77 | r_4_78 | r_4_79 | r_4_80 | r_4_81 | r_4_82 | r_4_83 | r_4_84 | r_4_85 | r_4_86 | r_4_87 | r_4_88 | r_4_89 | r_4_90 | r_4_91 | r_4_92 | r_4_93 | r_4_94 | r_4_95 | r_4_96 | r_4_97 | r_4_98 | r_4_99 | r_4_100, r_5_0 | r_5_1 | r_5_2 | r_5_3 | r_5_4 | r_5_5 | r_5_6 | r_5_7 | r_5_8 | r_5_9 | r_5_10 | r_5_11 | r_5_12 | r_5_13 | r_5_14 | r_5_15 | r_5_16 | r_5_17 | r_5_18 | r_5_19 | r_5_20 | r_5_21 | r_5_22 | r_5_23 | r_5_24 | r_5_25 | r_5_26 | r_5_27 | r_5_28 | r_5_29 | r_5_30 | r_5_31 | r_5_32 | r_5_33 | r_5_34 | r_5_35 | r_5_36 | r_5_37 | r_5_38 | r_5_39 | r_5_40 | r_5_41 | r_5_42 | r_5_43 | r_5_44 | r_5_45 | r_5_46 | r_5_47 | r_5_48 | r_5_49 | r_5_50 | r_5_51 | r_5_52 | r_5_53 | r_5_54 | r_5_55 | r_5_56 | r_5_57 | r_5_58 | r_5_59 | r_5_60 | r_5_61 | r_5_62 | r_5_63 | r_5_64 | r_5_65 | r_5_66 | r_5_67 | r_5_68 | r_5_69 | r_5_70 | r_5_71 | r_5_72 | r_5_73 | r_5_74 | r_5_75 | r_5_76 | r_5_77 | r_5_78 | r_5_79 | r_5_80 | r_5_81 | r_5_82 | r_5_83 | r_5_84 | r_5_85 | r_5_86 | r_5_87 | r_5_88 | r_5_89 | r_5_90 | r_5_91 | r_5_92 | r_5_93 | r_5_94 | r_5_95 | r_5_96 | r_5_97 | r_5_98 | r_5_99 | r_5_100};
  assign full_rank =  pivot_found == 6'b111111 ? 1'b1 : 1'b0;

  assign row0 = {r_0_0, r_0_1, r_0_2, r_0_3, r_0_4, r_0_5, r_0_6, r_0_7, r_0_8, r_0_9, r_0_10, r_0_11, r_0_12, r_0_13, r_0_14, r_0_15, r_0_16, r_0_17, r_0_18, r_0_19, r_0_20, r_0_21, r_0_22, r_0_23, r_0_24, r_0_25, r_0_26, r_0_27, r_0_28, r_0_29, r_0_30, r_0_31, r_0_32, r_0_33, r_0_34, r_0_35, r_0_36, r_0_37, r_0_38, r_0_39, r_0_40, r_0_41, r_0_42, r_0_43, r_0_44, r_0_45, r_0_46, r_0_47, r_0_48, r_0_49, r_0_50, r_0_51, r_0_52, r_0_53, r_0_54, r_0_55, r_0_56, r_0_57, r_0_58, r_0_59, r_0_60, r_0_61, r_0_62, r_0_63, r_0_64, r_0_65, r_0_66, r_0_67, r_0_68, r_0_69, r_0_70, r_0_71, r_0_72, r_0_73, r_0_74, r_0_75, r_0_76, r_0_77, r_0_78, r_0_79, r_0_80, r_0_81, r_0_82, r_0_83, r_0_84, r_0_85, r_0_86, r_0_87, r_0_88, r_0_89, r_0_90, r_0_91, r_0_92, r_0_93, r_0_94, r_0_95, r_0_96, r_0_97, r_0_98, r_0_99, r_0_100};
  assign row1 = {r_1_0, r_1_1, r_1_2, r_1_3, r_1_4, r_1_5, r_1_6, r_1_7, r_1_8, r_1_9, r_1_10, r_1_11, r_1_12, r_1_13, r_1_14, r_1_15, r_1_16, r_1_17, r_1_18, r_1_19, r_1_20, r_1_21, r_1_22, r_1_23, r_1_24, r_1_25, r_1_26, r_1_27, r_1_28, r_1_29, r_1_30, r_1_31, r_1_32, r_1_33, r_1_34, r_1_35, r_1_36, r_1_37, r_1_38, r_1_39, r_1_40, r_1_41, r_1_42, r_1_43, r_1_44, r_1_45, r_1_46, r_1_47, r_1_48, r_1_49, r_1_50, r_1_51, r_1_52, r_1_53, r_1_54, r_1_55, r_1_56, r_1_57, r_1_58, r_1_59, r_1_60, r_1_61, r_1_62, r_1_63, r_1_64, r_1_65, r_1_66, r_1_67, r_1_68, r_1_69, r_1_70, r_1_71, r_1_72, r_1_73, r_1_74, r_1_75, r_1_76, r_1_77, r_1_78, r_1_79, r_1_80, r_1_81, r_1_82, r_1_83, r_1_84, r_1_85, r_1_86, r_1_87, r_1_88, r_1_89, r_1_90, r_1_91, r_1_92, r_1_93, r_1_94, r_1_95, r_1_96, r_1_97, r_1_98, r_1_99, r_1_100};
  assign row2 = {r_2_0, r_2_1, r_2_2, r_2_3, r_2_4, r_2_5, r_2_6, r_2_7, r_2_8, r_2_9, r_2_10, r_2_11, r_2_12, r_2_13, r_2_14, r_2_15, r_2_16, r_2_17, r_2_18, r_2_19, r_2_20, r_2_21, r_2_22, r_2_23, r_2_24, r_2_25, r_2_26, r_2_27, r_2_28, r_2_29, r_2_30, r_2_31, r_2_32, r_2_33, r_2_34, r_2_35, r_2_36, r_2_37, r_2_38, r_2_39, r_2_40, r_2_41, r_2_42, r_2_43, r_2_44, r_2_45, r_2_46, r_2_47, r_2_48, r_2_49, r_2_50, r_2_51, r_2_52, r_2_53, r_2_54, r_2_55, r_2_56, r_2_57, r_2_58, r_2_59, r_2_60, r_2_61, r_2_62, r_2_63, r_2_64, r_2_65, r_2_66, r_2_67, r_2_68, r_2_69, r_2_70, r_2_71, r_2_72, r_2_73, r_2_74, r_2_75, r_2_76, r_2_77, r_2_78, r_2_79, r_2_80, r_2_81, r_2_82, r_2_83, r_2_84, r_2_85, r_2_86, r_2_87, r_2_88, r_2_89, r_2_90, r_2_91, r_2_92, r_2_93, r_2_94, r_2_95, r_2_96, r_2_97, r_2_98, r_2_99, r_2_100};
  assign row3 = {r_3_0, r_3_1, r_3_2, r_3_3, r_3_4, r_3_5, r_3_6, r_3_7, r_3_8, r_3_9, r_3_10, r_3_11, r_3_12, r_3_13, r_3_14, r_3_15, r_3_16, r_3_17, r_3_18, r_3_19, r_3_20, r_3_21, r_3_22, r_3_23, r_3_24, r_3_25, r_3_26, r_3_27, r_3_28, r_3_29, r_3_30, r_3_31, r_3_32, r_3_33, r_3_34, r_3_35, r_3_36, r_3_37, r_3_38, r_3_39, r_3_40, r_3_41, r_3_42, r_3_43, r_3_44, r_3_45, r_3_46, r_3_47, r_3_48, r_3_49, r_3_50, r_3_51, r_3_52, r_3_53, r_3_54, r_3_55, r_3_56, r_3_57, r_3_58, r_3_59, r_3_60, r_3_61, r_3_62, r_3_63, r_3_64, r_3_65, r_3_66, r_3_67, r_3_68, r_3_69, r_3_70, r_3_71, r_3_72, r_3_73, r_3_74, r_3_75, r_3_76, r_3_77, r_3_78, r_3_79, r_3_80, r_3_81, r_3_82, r_3_83, r_3_84, r_3_85, r_3_86, r_3_87, r_3_88, r_3_89, r_3_90, r_3_91, r_3_92, r_3_93, r_3_94, r_3_95, r_3_96, r_3_97, r_3_98, r_3_99, r_3_100};
  assign row4 = {r_4_0, r_4_1, r_4_2, r_4_3, r_4_4, r_4_5, r_4_6, r_4_7, r_4_8, r_4_9, r_4_10, r_4_11, r_4_12, r_4_13, r_4_14, r_4_15, r_4_16, r_4_17, r_4_18, r_4_19, r_4_20, r_4_21, r_4_22, r_4_23, r_4_24, r_4_25, r_4_26, r_4_27, r_4_28, r_4_29, r_4_30, r_4_31, r_4_32, r_4_33, r_4_34, r_4_35, r_4_36, r_4_37, r_4_38, r_4_39, r_4_40, r_4_41, r_4_42, r_4_43, r_4_44, r_4_45, r_4_46, r_4_47, r_4_48, r_4_49, r_4_50, r_4_51, r_4_52, r_4_53, r_4_54, r_4_55, r_4_56, r_4_57, r_4_58, r_4_59, r_4_60, r_4_61, r_4_62, r_4_63, r_4_64, r_4_65, r_4_66, r_4_67, r_4_68, r_4_69, r_4_70, r_4_71, r_4_72, r_4_73, r_4_74, r_4_75, r_4_76, r_4_77, r_4_78, r_4_79, r_4_80, r_4_81, r_4_82, r_4_83, r_4_84, r_4_85, r_4_86, r_4_87, r_4_88, r_4_89, r_4_90, r_4_91, r_4_92, r_4_93, r_4_94, r_4_95, r_4_96, r_4_97, r_4_98, r_4_99, r_4_100};
  assign row5 = {r_5_0, r_5_1, r_5_2, r_5_3, r_5_4, r_5_5, r_5_6, r_5_7, r_5_8, r_5_9, r_5_10, r_5_11, r_5_12, r_5_13, r_5_14, r_5_15, r_5_16, r_5_17, r_5_18, r_5_19, r_5_20, r_5_21, r_5_22, r_5_23, r_5_24, r_5_25, r_5_26, r_5_27, r_5_28, r_5_29, r_5_30, r_5_31, r_5_32, r_5_33, r_5_34, r_5_35, r_5_36, r_5_37, r_5_38, r_5_39, r_5_40, r_5_41, r_5_42, r_5_43, r_5_44, r_5_45, r_5_46, r_5_47, r_5_48, r_5_49, r_5_50, r_5_51, r_5_52, r_5_53, r_5_54, r_5_55, r_5_56, r_5_57, r_5_58, r_5_59, r_5_60, r_5_61, r_5_62, r_5_63, r_5_64, r_5_65, r_5_66, r_5_67, r_5_68, r_5_69, r_5_70, r_5_71, r_5_72, r_5_73, r_5_74, r_5_75, r_5_76, r_5_77, r_5_78, r_5_79, r_5_80, r_5_81, r_5_82, r_5_83, r_5_84, r_5_85, r_5_86, r_5_87, r_5_88, r_5_89, r_5_90, r_5_91, r_5_92, r_5_93, r_5_94, r_5_95, r_5_96, r_5_97, r_5_98, r_5_99, r_5_100};

  always @(posedge clk) begin
      finish <= ~mode ? start_out_5_100: start_out_0_99;
  end

   //output regular form from skewed form via pipelining
 reg [100:1] result_col0;
 reg [99:1] result_col1;
 reg [98:1] result_col2;
 reg [97:1] result_col3;
 reg [96:1] result_col4;
 reg [95:1] result_col5;
 reg [94:1] result_col6;
 reg [93:1] result_col7;
 reg [92:1] result_col8;
 reg [91:1] result_col9;
 reg [90:1] result_col10;
 reg [89:1] result_col11;
 reg [88:1] result_col12;
 reg [87:1] result_col13;
 reg [86:1] result_col14;
 reg [85:1] result_col15;
 reg [84:1] result_col16;
 reg [83:1] result_col17;
 reg [82:1] result_col18;
 reg [81:1] result_col19;
 reg [80:1] result_col20;
 reg [79:1] result_col21;
 reg [78:1] result_col22;
 reg [77:1] result_col23;
 reg [76:1] result_col24;
 reg [75:1] result_col25;
 reg [74:1] result_col26;
 reg [73:1] result_col27;
 reg [72:1] result_col28;
 reg [71:1] result_col29;
 reg [70:1] result_col30;
 reg [69:1] result_col31;
 reg [68:1] result_col32;
 reg [67:1] result_col33;
 reg [66:1] result_col34;
 reg [65:1] result_col35;
 reg [64:1] result_col36;
 reg [63:1] result_col37;
 reg [62:1] result_col38;
 reg [61:1] result_col39;
 reg [60:1] result_col40;
 reg [59:1] result_col41;
 reg [58:1] result_col42;
 reg [57:1] result_col43;
 reg [56:1] result_col44;
 reg [55:1] result_col45;
 reg [54:1] result_col46;
 reg [53:1] result_col47;
 reg [52:1] result_col48;
 reg [51:1] result_col49;
 reg [50:1] result_col50;
 reg [49:1] result_col51;
 reg [48:1] result_col52;
 reg [47:1] result_col53;
 reg [46:1] result_col54;
 reg [45:1] result_col55;
 reg [44:1] result_col56;
 reg [43:1] result_col57;
 reg [42:1] result_col58;
 reg [41:1] result_col59;
 reg [40:1] result_col60;
 reg [39:1] result_col61;
 reg [38:1] result_col62;
 reg [37:1] result_col63;
 reg [36:1] result_col64;
 reg [35:1] result_col65;
 reg [34:1] result_col66;
 reg [33:1] result_col67;
 reg [32:1] result_col68;
 reg [31:1] result_col69;
 reg [30:1] result_col70;
 reg [29:1] result_col71;
 reg [28:1] result_col72;
 reg [27:1] result_col73;
 reg [26:1] result_col74;
 reg [25:1] result_col75;
 reg [24:1] result_col76;
 reg [23:1] result_col77;
 reg [22:1] result_col78;
 reg [21:1] result_col79;
 reg [20:1] result_col80;
 reg [19:1] result_col81;
 reg [18:1] result_col82;
 reg [17:1] result_col83;
 reg [16:1] result_col84;
 reg [15:1] result_col85;
 reg [14:1] result_col86;
 reg [13:1] result_col87;
 reg [12:1] result_col88;
 reg [11:1] result_col89;
 reg [10:1] result_col90;
 reg [9:1] result_col91;
 reg [8:1] result_col92;
 reg [7:1] result_col93;
 reg [6:1] result_col94;
 reg [5:1] result_col95;
 reg [4:1] result_col96;
 reg [3:1] result_col97;
 reg [2:1] result_col98;
 reg [1:1] result_col99;
 wire result_col100;

 assign result_col100 = data_out_5_100;

  always @(posedge clk) begin
   result_col0[1] <= data_out_5_0;
   result_col0[2] <= result_col0[1];
   result_col0[3] <= result_col0[2];
   result_col0[4] <= result_col0[3];
   result_col0[5] <= result_col0[4];
   result_col0[6] <= result_col0[5];
   result_col0[7] <= result_col0[6];
   result_col0[8] <= result_col0[7];
   result_col0[9] <= result_col0[8];
   result_col0[10] <= result_col0[9];
   result_col0[11] <= result_col0[10];
   result_col0[12] <= result_col0[11];
   result_col0[13] <= result_col0[12];
   result_col0[14] <= result_col0[13];
   result_col0[15] <= result_col0[14];
   result_col0[16] <= result_col0[15];
   result_col0[17] <= result_col0[16];
   result_col0[18] <= result_col0[17];
   result_col0[19] <= result_col0[18];
   result_col0[20] <= result_col0[19];
   result_col0[21] <= result_col0[20];
   result_col0[22] <= result_col0[21];
   result_col0[23] <= result_col0[22];
   result_col0[24] <= result_col0[23];
   result_col0[25] <= result_col0[24];
   result_col0[26] <= result_col0[25];
   result_col0[27] <= result_col0[26];
   result_col0[28] <= result_col0[27];
   result_col0[29] <= result_col0[28];
   result_col0[30] <= result_col0[29];
   result_col0[31] <= result_col0[30];
   result_col0[32] <= result_col0[31];
   result_col0[33] <= result_col0[32];
   result_col0[34] <= result_col0[33];
   result_col0[35] <= result_col0[34];
   result_col0[36] <= result_col0[35];
   result_col0[37] <= result_col0[36];
   result_col0[38] <= result_col0[37];
   result_col0[39] <= result_col0[38];
   result_col0[40] <= result_col0[39];
   result_col0[41] <= result_col0[40];
   result_col0[42] <= result_col0[41];
   result_col0[43] <= result_col0[42];
   result_col0[44] <= result_col0[43];
   result_col0[45] <= result_col0[44];
   result_col0[46] <= result_col0[45];
   result_col0[47] <= result_col0[46];
   result_col0[48] <= result_col0[47];
   result_col0[49] <= result_col0[48];
   result_col0[50] <= result_col0[49];
   result_col0[51] <= result_col0[50];
   result_col0[52] <= result_col0[51];
   result_col0[53] <= result_col0[52];
   result_col0[54] <= result_col0[53];
   result_col0[55] <= result_col0[54];
   result_col0[56] <= result_col0[55];
   result_col0[57] <= result_col0[56];
   result_col0[58] <= result_col0[57];
   result_col0[59] <= result_col0[58];
   result_col0[60] <= result_col0[59];
   result_col0[61] <= result_col0[60];
   result_col0[62] <= result_col0[61];
   result_col0[63] <= result_col0[62];
   result_col0[64] <= result_col0[63];
   result_col0[65] <= result_col0[64];
   result_col0[66] <= result_col0[65];
   result_col0[67] <= result_col0[66];
   result_col0[68] <= result_col0[67];
   result_col0[69] <= result_col0[68];
   result_col0[70] <= result_col0[69];
   result_col0[71] <= result_col0[70];
   result_col0[72] <= result_col0[71];
   result_col0[73] <= result_col0[72];
   result_col0[74] <= result_col0[73];
   result_col0[75] <= result_col0[74];
   result_col0[76] <= result_col0[75];
   result_col0[77] <= result_col0[76];
   result_col0[78] <= result_col0[77];
   result_col0[79] <= result_col0[78];
   result_col0[80] <= result_col0[79];
   result_col0[81] <= result_col0[80];
   result_col0[82] <= result_col0[81];
   result_col0[83] <= result_col0[82];
   result_col0[84] <= result_col0[83];
   result_col0[85] <= result_col0[84];
   result_col0[86] <= result_col0[85];
   result_col0[87] <= result_col0[86];
   result_col0[88] <= result_col0[87];
   result_col0[89] <= result_col0[88];
   result_col0[90] <= result_col0[89];
   result_col0[91] <= result_col0[90];
   result_col0[92] <= result_col0[91];
   result_col0[93] <= result_col0[92];
   result_col0[94] <= result_col0[93];
   result_col0[95] <= result_col0[94];
   result_col0[96] <= result_col0[95];
   result_col0[97] <= result_col0[96];
   result_col0[98] <= result_col0[97];
   result_col0[99] <= result_col0[98];
   result_col0[100] <= result_col0[99];

   result_col1[1] <= data_out_5_1;
   result_col1[2] <= result_col1[1];
   result_col1[3] <= result_col1[2];
   result_col1[4] <= result_col1[3];
   result_col1[5] <= result_col1[4];
   result_col1[6] <= result_col1[5];
   result_col1[7] <= result_col1[6];
   result_col1[8] <= result_col1[7];
   result_col1[9] <= result_col1[8];
   result_col1[10] <= result_col1[9];
   result_col1[11] <= result_col1[10];
   result_col1[12] <= result_col1[11];
   result_col1[13] <= result_col1[12];
   result_col1[14] <= result_col1[13];
   result_col1[15] <= result_col1[14];
   result_col1[16] <= result_col1[15];
   result_col1[17] <= result_col1[16];
   result_col1[18] <= result_col1[17];
   result_col1[19] <= result_col1[18];
   result_col1[20] <= result_col1[19];
   result_col1[21] <= result_col1[20];
   result_col1[22] <= result_col1[21];
   result_col1[23] <= result_col1[22];
   result_col1[24] <= result_col1[23];
   result_col1[25] <= result_col1[24];
   result_col1[26] <= result_col1[25];
   result_col1[27] <= result_col1[26];
   result_col1[28] <= result_col1[27];
   result_col1[29] <= result_col1[28];
   result_col1[30] <= result_col1[29];
   result_col1[31] <= result_col1[30];
   result_col1[32] <= result_col1[31];
   result_col1[33] <= result_col1[32];
   result_col1[34] <= result_col1[33];
   result_col1[35] <= result_col1[34];
   result_col1[36] <= result_col1[35];
   result_col1[37] <= result_col1[36];
   result_col1[38] <= result_col1[37];
   result_col1[39] <= result_col1[38];
   result_col1[40] <= result_col1[39];
   result_col1[41] <= result_col1[40];
   result_col1[42] <= result_col1[41];
   result_col1[43] <= result_col1[42];
   result_col1[44] <= result_col1[43];
   result_col1[45] <= result_col1[44];
   result_col1[46] <= result_col1[45];
   result_col1[47] <= result_col1[46];
   result_col1[48] <= result_col1[47];
   result_col1[49] <= result_col1[48];
   result_col1[50] <= result_col1[49];
   result_col1[51] <= result_col1[50];
   result_col1[52] <= result_col1[51];
   result_col1[53] <= result_col1[52];
   result_col1[54] <= result_col1[53];
   result_col1[55] <= result_col1[54];
   result_col1[56] <= result_col1[55];
   result_col1[57] <= result_col1[56];
   result_col1[58] <= result_col1[57];
   result_col1[59] <= result_col1[58];
   result_col1[60] <= result_col1[59];
   result_col1[61] <= result_col1[60];
   result_col1[62] <= result_col1[61];
   result_col1[63] <= result_col1[62];
   result_col1[64] <= result_col1[63];
   result_col1[65] <= result_col1[64];
   result_col1[66] <= result_col1[65];
   result_col1[67] <= result_col1[66];
   result_col1[68] <= result_col1[67];
   result_col1[69] <= result_col1[68];
   result_col1[70] <= result_col1[69];
   result_col1[71] <= result_col1[70];
   result_col1[72] <= result_col1[71];
   result_col1[73] <= result_col1[72];
   result_col1[74] <= result_col1[73];
   result_col1[75] <= result_col1[74];
   result_col1[76] <= result_col1[75];
   result_col1[77] <= result_col1[76];
   result_col1[78] <= result_col1[77];
   result_col1[79] <= result_col1[78];
   result_col1[80] <= result_col1[79];
   result_col1[81] <= result_col1[80];
   result_col1[82] <= result_col1[81];
   result_col1[83] <= result_col1[82];
   result_col1[84] <= result_col1[83];
   result_col1[85] <= result_col1[84];
   result_col1[86] <= result_col1[85];
   result_col1[87] <= result_col1[86];
   result_col1[88] <= result_col1[87];
   result_col1[89] <= result_col1[88];
   result_col1[90] <= result_col1[89];
   result_col1[91] <= result_col1[90];
   result_col1[92] <= result_col1[91];
   result_col1[93] <= result_col1[92];
   result_col1[94] <= result_col1[93];
   result_col1[95] <= result_col1[94];
   result_col1[96] <= result_col1[95];
   result_col1[97] <= result_col1[96];
   result_col1[98] <= result_col1[97];
   result_col1[99] <= result_col1[98];

   result_col2[1] <= data_out_5_2;
   result_col2[2] <= result_col2[1];
   result_col2[3] <= result_col2[2];
   result_col2[4] <= result_col2[3];
   result_col2[5] <= result_col2[4];
   result_col2[6] <= result_col2[5];
   result_col2[7] <= result_col2[6];
   result_col2[8] <= result_col2[7];
   result_col2[9] <= result_col2[8];
   result_col2[10] <= result_col2[9];
   result_col2[11] <= result_col2[10];
   result_col2[12] <= result_col2[11];
   result_col2[13] <= result_col2[12];
   result_col2[14] <= result_col2[13];
   result_col2[15] <= result_col2[14];
   result_col2[16] <= result_col2[15];
   result_col2[17] <= result_col2[16];
   result_col2[18] <= result_col2[17];
   result_col2[19] <= result_col2[18];
   result_col2[20] <= result_col2[19];
   result_col2[21] <= result_col2[20];
   result_col2[22] <= result_col2[21];
   result_col2[23] <= result_col2[22];
   result_col2[24] <= result_col2[23];
   result_col2[25] <= result_col2[24];
   result_col2[26] <= result_col2[25];
   result_col2[27] <= result_col2[26];
   result_col2[28] <= result_col2[27];
   result_col2[29] <= result_col2[28];
   result_col2[30] <= result_col2[29];
   result_col2[31] <= result_col2[30];
   result_col2[32] <= result_col2[31];
   result_col2[33] <= result_col2[32];
   result_col2[34] <= result_col2[33];
   result_col2[35] <= result_col2[34];
   result_col2[36] <= result_col2[35];
   result_col2[37] <= result_col2[36];
   result_col2[38] <= result_col2[37];
   result_col2[39] <= result_col2[38];
   result_col2[40] <= result_col2[39];
   result_col2[41] <= result_col2[40];
   result_col2[42] <= result_col2[41];
   result_col2[43] <= result_col2[42];
   result_col2[44] <= result_col2[43];
   result_col2[45] <= result_col2[44];
   result_col2[46] <= result_col2[45];
   result_col2[47] <= result_col2[46];
   result_col2[48] <= result_col2[47];
   result_col2[49] <= result_col2[48];
   result_col2[50] <= result_col2[49];
   result_col2[51] <= result_col2[50];
   result_col2[52] <= result_col2[51];
   result_col2[53] <= result_col2[52];
   result_col2[54] <= result_col2[53];
   result_col2[55] <= result_col2[54];
   result_col2[56] <= result_col2[55];
   result_col2[57] <= result_col2[56];
   result_col2[58] <= result_col2[57];
   result_col2[59] <= result_col2[58];
   result_col2[60] <= result_col2[59];
   result_col2[61] <= result_col2[60];
   result_col2[62] <= result_col2[61];
   result_col2[63] <= result_col2[62];
   result_col2[64] <= result_col2[63];
   result_col2[65] <= result_col2[64];
   result_col2[66] <= result_col2[65];
   result_col2[67] <= result_col2[66];
   result_col2[68] <= result_col2[67];
   result_col2[69] <= result_col2[68];
   result_col2[70] <= result_col2[69];
   result_col2[71] <= result_col2[70];
   result_col2[72] <= result_col2[71];
   result_col2[73] <= result_col2[72];
   result_col2[74] <= result_col2[73];
   result_col2[75] <= result_col2[74];
   result_col2[76] <= result_col2[75];
   result_col2[77] <= result_col2[76];
   result_col2[78] <= result_col2[77];
   result_col2[79] <= result_col2[78];
   result_col2[80] <= result_col2[79];
   result_col2[81] <= result_col2[80];
   result_col2[82] <= result_col2[81];
   result_col2[83] <= result_col2[82];
   result_col2[84] <= result_col2[83];
   result_col2[85] <= result_col2[84];
   result_col2[86] <= result_col2[85];
   result_col2[87] <= result_col2[86];
   result_col2[88] <= result_col2[87];
   result_col2[89] <= result_col2[88];
   result_col2[90] <= result_col2[89];
   result_col2[91] <= result_col2[90];
   result_col2[92] <= result_col2[91];
   result_col2[93] <= result_col2[92];
   result_col2[94] <= result_col2[93];
   result_col2[95] <= result_col2[94];
   result_col2[96] <= result_col2[95];
   result_col2[97] <= result_col2[96];
   result_col2[98] <= result_col2[97];

   result_col3[1] <= data_out_5_3;
   result_col3[2] <= result_col3[1];
   result_col3[3] <= result_col3[2];
   result_col3[4] <= result_col3[3];
   result_col3[5] <= result_col3[4];
   result_col3[6] <= result_col3[5];
   result_col3[7] <= result_col3[6];
   result_col3[8] <= result_col3[7];
   result_col3[9] <= result_col3[8];
   result_col3[10] <= result_col3[9];
   result_col3[11] <= result_col3[10];
   result_col3[12] <= result_col3[11];
   result_col3[13] <= result_col3[12];
   result_col3[14] <= result_col3[13];
   result_col3[15] <= result_col3[14];
   result_col3[16] <= result_col3[15];
   result_col3[17] <= result_col3[16];
   result_col3[18] <= result_col3[17];
   result_col3[19] <= result_col3[18];
   result_col3[20] <= result_col3[19];
   result_col3[21] <= result_col3[20];
   result_col3[22] <= result_col3[21];
   result_col3[23] <= result_col3[22];
   result_col3[24] <= result_col3[23];
   result_col3[25] <= result_col3[24];
   result_col3[26] <= result_col3[25];
   result_col3[27] <= result_col3[26];
   result_col3[28] <= result_col3[27];
   result_col3[29] <= result_col3[28];
   result_col3[30] <= result_col3[29];
   result_col3[31] <= result_col3[30];
   result_col3[32] <= result_col3[31];
   result_col3[33] <= result_col3[32];
   result_col3[34] <= result_col3[33];
   result_col3[35] <= result_col3[34];
   result_col3[36] <= result_col3[35];
   result_col3[37] <= result_col3[36];
   result_col3[38] <= result_col3[37];
   result_col3[39] <= result_col3[38];
   result_col3[40] <= result_col3[39];
   result_col3[41] <= result_col3[40];
   result_col3[42] <= result_col3[41];
   result_col3[43] <= result_col3[42];
   result_col3[44] <= result_col3[43];
   result_col3[45] <= result_col3[44];
   result_col3[46] <= result_col3[45];
   result_col3[47] <= result_col3[46];
   result_col3[48] <= result_col3[47];
   result_col3[49] <= result_col3[48];
   result_col3[50] <= result_col3[49];
   result_col3[51] <= result_col3[50];
   result_col3[52] <= result_col3[51];
   result_col3[53] <= result_col3[52];
   result_col3[54] <= result_col3[53];
   result_col3[55] <= result_col3[54];
   result_col3[56] <= result_col3[55];
   result_col3[57] <= result_col3[56];
   result_col3[58] <= result_col3[57];
   result_col3[59] <= result_col3[58];
   result_col3[60] <= result_col3[59];
   result_col3[61] <= result_col3[60];
   result_col3[62] <= result_col3[61];
   result_col3[63] <= result_col3[62];
   result_col3[64] <= result_col3[63];
   result_col3[65] <= result_col3[64];
   result_col3[66] <= result_col3[65];
   result_col3[67] <= result_col3[66];
   result_col3[68] <= result_col3[67];
   result_col3[69] <= result_col3[68];
   result_col3[70] <= result_col3[69];
   result_col3[71] <= result_col3[70];
   result_col3[72] <= result_col3[71];
   result_col3[73] <= result_col3[72];
   result_col3[74] <= result_col3[73];
   result_col3[75] <= result_col3[74];
   result_col3[76] <= result_col3[75];
   result_col3[77] <= result_col3[76];
   result_col3[78] <= result_col3[77];
   result_col3[79] <= result_col3[78];
   result_col3[80] <= result_col3[79];
   result_col3[81] <= result_col3[80];
   result_col3[82] <= result_col3[81];
   result_col3[83] <= result_col3[82];
   result_col3[84] <= result_col3[83];
   result_col3[85] <= result_col3[84];
   result_col3[86] <= result_col3[85];
   result_col3[87] <= result_col3[86];
   result_col3[88] <= result_col3[87];
   result_col3[89] <= result_col3[88];
   result_col3[90] <= result_col3[89];
   result_col3[91] <= result_col3[90];
   result_col3[92] <= result_col3[91];
   result_col3[93] <= result_col3[92];
   result_col3[94] <= result_col3[93];
   result_col3[95] <= result_col3[94];
   result_col3[96] <= result_col3[95];
   result_col3[97] <= result_col3[96];

   result_col4[1] <= data_out_5_4;
   result_col4[2] <= result_col4[1];
   result_col4[3] <= result_col4[2];
   result_col4[4] <= result_col4[3];
   result_col4[5] <= result_col4[4];
   result_col4[6] <= result_col4[5];
   result_col4[7] <= result_col4[6];
   result_col4[8] <= result_col4[7];
   result_col4[9] <= result_col4[8];
   result_col4[10] <= result_col4[9];
   result_col4[11] <= result_col4[10];
   result_col4[12] <= result_col4[11];
   result_col4[13] <= result_col4[12];
   result_col4[14] <= result_col4[13];
   result_col4[15] <= result_col4[14];
   result_col4[16] <= result_col4[15];
   result_col4[17] <= result_col4[16];
   result_col4[18] <= result_col4[17];
   result_col4[19] <= result_col4[18];
   result_col4[20] <= result_col4[19];
   result_col4[21] <= result_col4[20];
   result_col4[22] <= result_col4[21];
   result_col4[23] <= result_col4[22];
   result_col4[24] <= result_col4[23];
   result_col4[25] <= result_col4[24];
   result_col4[26] <= result_col4[25];
   result_col4[27] <= result_col4[26];
   result_col4[28] <= result_col4[27];
   result_col4[29] <= result_col4[28];
   result_col4[30] <= result_col4[29];
   result_col4[31] <= result_col4[30];
   result_col4[32] <= result_col4[31];
   result_col4[33] <= result_col4[32];
   result_col4[34] <= result_col4[33];
   result_col4[35] <= result_col4[34];
   result_col4[36] <= result_col4[35];
   result_col4[37] <= result_col4[36];
   result_col4[38] <= result_col4[37];
   result_col4[39] <= result_col4[38];
   result_col4[40] <= result_col4[39];
   result_col4[41] <= result_col4[40];
   result_col4[42] <= result_col4[41];
   result_col4[43] <= result_col4[42];
   result_col4[44] <= result_col4[43];
   result_col4[45] <= result_col4[44];
   result_col4[46] <= result_col4[45];
   result_col4[47] <= result_col4[46];
   result_col4[48] <= result_col4[47];
   result_col4[49] <= result_col4[48];
   result_col4[50] <= result_col4[49];
   result_col4[51] <= result_col4[50];
   result_col4[52] <= result_col4[51];
   result_col4[53] <= result_col4[52];
   result_col4[54] <= result_col4[53];
   result_col4[55] <= result_col4[54];
   result_col4[56] <= result_col4[55];
   result_col4[57] <= result_col4[56];
   result_col4[58] <= result_col4[57];
   result_col4[59] <= result_col4[58];
   result_col4[60] <= result_col4[59];
   result_col4[61] <= result_col4[60];
   result_col4[62] <= result_col4[61];
   result_col4[63] <= result_col4[62];
   result_col4[64] <= result_col4[63];
   result_col4[65] <= result_col4[64];
   result_col4[66] <= result_col4[65];
   result_col4[67] <= result_col4[66];
   result_col4[68] <= result_col4[67];
   result_col4[69] <= result_col4[68];
   result_col4[70] <= result_col4[69];
   result_col4[71] <= result_col4[70];
   result_col4[72] <= result_col4[71];
   result_col4[73] <= result_col4[72];
   result_col4[74] <= result_col4[73];
   result_col4[75] <= result_col4[74];
   result_col4[76] <= result_col4[75];
   result_col4[77] <= result_col4[76];
   result_col4[78] <= result_col4[77];
   result_col4[79] <= result_col4[78];
   result_col4[80] <= result_col4[79];
   result_col4[81] <= result_col4[80];
   result_col4[82] <= result_col4[81];
   result_col4[83] <= result_col4[82];
   result_col4[84] <= result_col4[83];
   result_col4[85] <= result_col4[84];
   result_col4[86] <= result_col4[85];
   result_col4[87] <= result_col4[86];
   result_col4[88] <= result_col4[87];
   result_col4[89] <= result_col4[88];
   result_col4[90] <= result_col4[89];
   result_col4[91] <= result_col4[90];
   result_col4[92] <= result_col4[91];
   result_col4[93] <= result_col4[92];
   result_col4[94] <= result_col4[93];
   result_col4[95] <= result_col4[94];
   result_col4[96] <= result_col4[95];

   result_col5[1] <= data_out_5_5;
   result_col5[2] <= result_col5[1];
   result_col5[3] <= result_col5[2];
   result_col5[4] <= result_col5[3];
   result_col5[5] <= result_col5[4];
   result_col5[6] <= result_col5[5];
   result_col5[7] <= result_col5[6];
   result_col5[8] <= result_col5[7];
   result_col5[9] <= result_col5[8];
   result_col5[10] <= result_col5[9];
   result_col5[11] <= result_col5[10];
   result_col5[12] <= result_col5[11];
   result_col5[13] <= result_col5[12];
   result_col5[14] <= result_col5[13];
   result_col5[15] <= result_col5[14];
   result_col5[16] <= result_col5[15];
   result_col5[17] <= result_col5[16];
   result_col5[18] <= result_col5[17];
   result_col5[19] <= result_col5[18];
   result_col5[20] <= result_col5[19];
   result_col5[21] <= result_col5[20];
   result_col5[22] <= result_col5[21];
   result_col5[23] <= result_col5[22];
   result_col5[24] <= result_col5[23];
   result_col5[25] <= result_col5[24];
   result_col5[26] <= result_col5[25];
   result_col5[27] <= result_col5[26];
   result_col5[28] <= result_col5[27];
   result_col5[29] <= result_col5[28];
   result_col5[30] <= result_col5[29];
   result_col5[31] <= result_col5[30];
   result_col5[32] <= result_col5[31];
   result_col5[33] <= result_col5[32];
   result_col5[34] <= result_col5[33];
   result_col5[35] <= result_col5[34];
   result_col5[36] <= result_col5[35];
   result_col5[37] <= result_col5[36];
   result_col5[38] <= result_col5[37];
   result_col5[39] <= result_col5[38];
   result_col5[40] <= result_col5[39];
   result_col5[41] <= result_col5[40];
   result_col5[42] <= result_col5[41];
   result_col5[43] <= result_col5[42];
   result_col5[44] <= result_col5[43];
   result_col5[45] <= result_col5[44];
   result_col5[46] <= result_col5[45];
   result_col5[47] <= result_col5[46];
   result_col5[48] <= result_col5[47];
   result_col5[49] <= result_col5[48];
   result_col5[50] <= result_col5[49];
   result_col5[51] <= result_col5[50];
   result_col5[52] <= result_col5[51];
   result_col5[53] <= result_col5[52];
   result_col5[54] <= result_col5[53];
   result_col5[55] <= result_col5[54];
   result_col5[56] <= result_col5[55];
   result_col5[57] <= result_col5[56];
   result_col5[58] <= result_col5[57];
   result_col5[59] <= result_col5[58];
   result_col5[60] <= result_col5[59];
   result_col5[61] <= result_col5[60];
   result_col5[62] <= result_col5[61];
   result_col5[63] <= result_col5[62];
   result_col5[64] <= result_col5[63];
   result_col5[65] <= result_col5[64];
   result_col5[66] <= result_col5[65];
   result_col5[67] <= result_col5[66];
   result_col5[68] <= result_col5[67];
   result_col5[69] <= result_col5[68];
   result_col5[70] <= result_col5[69];
   result_col5[71] <= result_col5[70];
   result_col5[72] <= result_col5[71];
   result_col5[73] <= result_col5[72];
   result_col5[74] <= result_col5[73];
   result_col5[75] <= result_col5[74];
   result_col5[76] <= result_col5[75];
   result_col5[77] <= result_col5[76];
   result_col5[78] <= result_col5[77];
   result_col5[79] <= result_col5[78];
   result_col5[80] <= result_col5[79];
   result_col5[81] <= result_col5[80];
   result_col5[82] <= result_col5[81];
   result_col5[83] <= result_col5[82];
   result_col5[84] <= result_col5[83];
   result_col5[85] <= result_col5[84];
   result_col5[86] <= result_col5[85];
   result_col5[87] <= result_col5[86];
   result_col5[88] <= result_col5[87];
   result_col5[89] <= result_col5[88];
   result_col5[90] <= result_col5[89];
   result_col5[91] <= result_col5[90];
   result_col5[92] <= result_col5[91];
   result_col5[93] <= result_col5[92];
   result_col5[94] <= result_col5[93];
   result_col5[95] <= result_col5[94];

   result_col6[1] <= data_out_5_6;
   result_col6[2] <= result_col6[1];
   result_col6[3] <= result_col6[2];
   result_col6[4] <= result_col6[3];
   result_col6[5] <= result_col6[4];
   result_col6[6] <= result_col6[5];
   result_col6[7] <= result_col6[6];
   result_col6[8] <= result_col6[7];
   result_col6[9] <= result_col6[8];
   result_col6[10] <= result_col6[9];
   result_col6[11] <= result_col6[10];
   result_col6[12] <= result_col6[11];
   result_col6[13] <= result_col6[12];
   result_col6[14] <= result_col6[13];
   result_col6[15] <= result_col6[14];
   result_col6[16] <= result_col6[15];
   result_col6[17] <= result_col6[16];
   result_col6[18] <= result_col6[17];
   result_col6[19] <= result_col6[18];
   result_col6[20] <= result_col6[19];
   result_col6[21] <= result_col6[20];
   result_col6[22] <= result_col6[21];
   result_col6[23] <= result_col6[22];
   result_col6[24] <= result_col6[23];
   result_col6[25] <= result_col6[24];
   result_col6[26] <= result_col6[25];
   result_col6[27] <= result_col6[26];
   result_col6[28] <= result_col6[27];
   result_col6[29] <= result_col6[28];
   result_col6[30] <= result_col6[29];
   result_col6[31] <= result_col6[30];
   result_col6[32] <= result_col6[31];
   result_col6[33] <= result_col6[32];
   result_col6[34] <= result_col6[33];
   result_col6[35] <= result_col6[34];
   result_col6[36] <= result_col6[35];
   result_col6[37] <= result_col6[36];
   result_col6[38] <= result_col6[37];
   result_col6[39] <= result_col6[38];
   result_col6[40] <= result_col6[39];
   result_col6[41] <= result_col6[40];
   result_col6[42] <= result_col6[41];
   result_col6[43] <= result_col6[42];
   result_col6[44] <= result_col6[43];
   result_col6[45] <= result_col6[44];
   result_col6[46] <= result_col6[45];
   result_col6[47] <= result_col6[46];
   result_col6[48] <= result_col6[47];
   result_col6[49] <= result_col6[48];
   result_col6[50] <= result_col6[49];
   result_col6[51] <= result_col6[50];
   result_col6[52] <= result_col6[51];
   result_col6[53] <= result_col6[52];
   result_col6[54] <= result_col6[53];
   result_col6[55] <= result_col6[54];
   result_col6[56] <= result_col6[55];
   result_col6[57] <= result_col6[56];
   result_col6[58] <= result_col6[57];
   result_col6[59] <= result_col6[58];
   result_col6[60] <= result_col6[59];
   result_col6[61] <= result_col6[60];
   result_col6[62] <= result_col6[61];
   result_col6[63] <= result_col6[62];
   result_col6[64] <= result_col6[63];
   result_col6[65] <= result_col6[64];
   result_col6[66] <= result_col6[65];
   result_col6[67] <= result_col6[66];
   result_col6[68] <= result_col6[67];
   result_col6[69] <= result_col6[68];
   result_col6[70] <= result_col6[69];
   result_col6[71] <= result_col6[70];
   result_col6[72] <= result_col6[71];
   result_col6[73] <= result_col6[72];
   result_col6[74] <= result_col6[73];
   result_col6[75] <= result_col6[74];
   result_col6[76] <= result_col6[75];
   result_col6[77] <= result_col6[76];
   result_col6[78] <= result_col6[77];
   result_col6[79] <= result_col6[78];
   result_col6[80] <= result_col6[79];
   result_col6[81] <= result_col6[80];
   result_col6[82] <= result_col6[81];
   result_col6[83] <= result_col6[82];
   result_col6[84] <= result_col6[83];
   result_col6[85] <= result_col6[84];
   result_col6[86] <= result_col6[85];
   result_col6[87] <= result_col6[86];
   result_col6[88] <= result_col6[87];
   result_col6[89] <= result_col6[88];
   result_col6[90] <= result_col6[89];
   result_col6[91] <= result_col6[90];
   result_col6[92] <= result_col6[91];
   result_col6[93] <= result_col6[92];
   result_col6[94] <= result_col6[93];

   result_col7[1] <= data_out_5_7;
   result_col7[2] <= result_col7[1];
   result_col7[3] <= result_col7[2];
   result_col7[4] <= result_col7[3];
   result_col7[5] <= result_col7[4];
   result_col7[6] <= result_col7[5];
   result_col7[7] <= result_col7[6];
   result_col7[8] <= result_col7[7];
   result_col7[9] <= result_col7[8];
   result_col7[10] <= result_col7[9];
   result_col7[11] <= result_col7[10];
   result_col7[12] <= result_col7[11];
   result_col7[13] <= result_col7[12];
   result_col7[14] <= result_col7[13];
   result_col7[15] <= result_col7[14];
   result_col7[16] <= result_col7[15];
   result_col7[17] <= result_col7[16];
   result_col7[18] <= result_col7[17];
   result_col7[19] <= result_col7[18];
   result_col7[20] <= result_col7[19];
   result_col7[21] <= result_col7[20];
   result_col7[22] <= result_col7[21];
   result_col7[23] <= result_col7[22];
   result_col7[24] <= result_col7[23];
   result_col7[25] <= result_col7[24];
   result_col7[26] <= result_col7[25];
   result_col7[27] <= result_col7[26];
   result_col7[28] <= result_col7[27];
   result_col7[29] <= result_col7[28];
   result_col7[30] <= result_col7[29];
   result_col7[31] <= result_col7[30];
   result_col7[32] <= result_col7[31];
   result_col7[33] <= result_col7[32];
   result_col7[34] <= result_col7[33];
   result_col7[35] <= result_col7[34];
   result_col7[36] <= result_col7[35];
   result_col7[37] <= result_col7[36];
   result_col7[38] <= result_col7[37];
   result_col7[39] <= result_col7[38];
   result_col7[40] <= result_col7[39];
   result_col7[41] <= result_col7[40];
   result_col7[42] <= result_col7[41];
   result_col7[43] <= result_col7[42];
   result_col7[44] <= result_col7[43];
   result_col7[45] <= result_col7[44];
   result_col7[46] <= result_col7[45];
   result_col7[47] <= result_col7[46];
   result_col7[48] <= result_col7[47];
   result_col7[49] <= result_col7[48];
   result_col7[50] <= result_col7[49];
   result_col7[51] <= result_col7[50];
   result_col7[52] <= result_col7[51];
   result_col7[53] <= result_col7[52];
   result_col7[54] <= result_col7[53];
   result_col7[55] <= result_col7[54];
   result_col7[56] <= result_col7[55];
   result_col7[57] <= result_col7[56];
   result_col7[58] <= result_col7[57];
   result_col7[59] <= result_col7[58];
   result_col7[60] <= result_col7[59];
   result_col7[61] <= result_col7[60];
   result_col7[62] <= result_col7[61];
   result_col7[63] <= result_col7[62];
   result_col7[64] <= result_col7[63];
   result_col7[65] <= result_col7[64];
   result_col7[66] <= result_col7[65];
   result_col7[67] <= result_col7[66];
   result_col7[68] <= result_col7[67];
   result_col7[69] <= result_col7[68];
   result_col7[70] <= result_col7[69];
   result_col7[71] <= result_col7[70];
   result_col7[72] <= result_col7[71];
   result_col7[73] <= result_col7[72];
   result_col7[74] <= result_col7[73];
   result_col7[75] <= result_col7[74];
   result_col7[76] <= result_col7[75];
   result_col7[77] <= result_col7[76];
   result_col7[78] <= result_col7[77];
   result_col7[79] <= result_col7[78];
   result_col7[80] <= result_col7[79];
   result_col7[81] <= result_col7[80];
   result_col7[82] <= result_col7[81];
   result_col7[83] <= result_col7[82];
   result_col7[84] <= result_col7[83];
   result_col7[85] <= result_col7[84];
   result_col7[86] <= result_col7[85];
   result_col7[87] <= result_col7[86];
   result_col7[88] <= result_col7[87];
   result_col7[89] <= result_col7[88];
   result_col7[90] <= result_col7[89];
   result_col7[91] <= result_col7[90];
   result_col7[92] <= result_col7[91];
   result_col7[93] <= result_col7[92];

   result_col8[1] <= data_out_5_8;
   result_col8[2] <= result_col8[1];
   result_col8[3] <= result_col8[2];
   result_col8[4] <= result_col8[3];
   result_col8[5] <= result_col8[4];
   result_col8[6] <= result_col8[5];
   result_col8[7] <= result_col8[6];
   result_col8[8] <= result_col8[7];
   result_col8[9] <= result_col8[8];
   result_col8[10] <= result_col8[9];
   result_col8[11] <= result_col8[10];
   result_col8[12] <= result_col8[11];
   result_col8[13] <= result_col8[12];
   result_col8[14] <= result_col8[13];
   result_col8[15] <= result_col8[14];
   result_col8[16] <= result_col8[15];
   result_col8[17] <= result_col8[16];
   result_col8[18] <= result_col8[17];
   result_col8[19] <= result_col8[18];
   result_col8[20] <= result_col8[19];
   result_col8[21] <= result_col8[20];
   result_col8[22] <= result_col8[21];
   result_col8[23] <= result_col8[22];
   result_col8[24] <= result_col8[23];
   result_col8[25] <= result_col8[24];
   result_col8[26] <= result_col8[25];
   result_col8[27] <= result_col8[26];
   result_col8[28] <= result_col8[27];
   result_col8[29] <= result_col8[28];
   result_col8[30] <= result_col8[29];
   result_col8[31] <= result_col8[30];
   result_col8[32] <= result_col8[31];
   result_col8[33] <= result_col8[32];
   result_col8[34] <= result_col8[33];
   result_col8[35] <= result_col8[34];
   result_col8[36] <= result_col8[35];
   result_col8[37] <= result_col8[36];
   result_col8[38] <= result_col8[37];
   result_col8[39] <= result_col8[38];
   result_col8[40] <= result_col8[39];
   result_col8[41] <= result_col8[40];
   result_col8[42] <= result_col8[41];
   result_col8[43] <= result_col8[42];
   result_col8[44] <= result_col8[43];
   result_col8[45] <= result_col8[44];
   result_col8[46] <= result_col8[45];
   result_col8[47] <= result_col8[46];
   result_col8[48] <= result_col8[47];
   result_col8[49] <= result_col8[48];
   result_col8[50] <= result_col8[49];
   result_col8[51] <= result_col8[50];
   result_col8[52] <= result_col8[51];
   result_col8[53] <= result_col8[52];
   result_col8[54] <= result_col8[53];
   result_col8[55] <= result_col8[54];
   result_col8[56] <= result_col8[55];
   result_col8[57] <= result_col8[56];
   result_col8[58] <= result_col8[57];
   result_col8[59] <= result_col8[58];
   result_col8[60] <= result_col8[59];
   result_col8[61] <= result_col8[60];
   result_col8[62] <= result_col8[61];
   result_col8[63] <= result_col8[62];
   result_col8[64] <= result_col8[63];
   result_col8[65] <= result_col8[64];
   result_col8[66] <= result_col8[65];
   result_col8[67] <= result_col8[66];
   result_col8[68] <= result_col8[67];
   result_col8[69] <= result_col8[68];
   result_col8[70] <= result_col8[69];
   result_col8[71] <= result_col8[70];
   result_col8[72] <= result_col8[71];
   result_col8[73] <= result_col8[72];
   result_col8[74] <= result_col8[73];
   result_col8[75] <= result_col8[74];
   result_col8[76] <= result_col8[75];
   result_col8[77] <= result_col8[76];
   result_col8[78] <= result_col8[77];
   result_col8[79] <= result_col8[78];
   result_col8[80] <= result_col8[79];
   result_col8[81] <= result_col8[80];
   result_col8[82] <= result_col8[81];
   result_col8[83] <= result_col8[82];
   result_col8[84] <= result_col8[83];
   result_col8[85] <= result_col8[84];
   result_col8[86] <= result_col8[85];
   result_col8[87] <= result_col8[86];
   result_col8[88] <= result_col8[87];
   result_col8[89] <= result_col8[88];
   result_col8[90] <= result_col8[89];
   result_col8[91] <= result_col8[90];
   result_col8[92] <= result_col8[91];

   result_col9[1] <= data_out_5_9;
   result_col9[2] <= result_col9[1];
   result_col9[3] <= result_col9[2];
   result_col9[4] <= result_col9[3];
   result_col9[5] <= result_col9[4];
   result_col9[6] <= result_col9[5];
   result_col9[7] <= result_col9[6];
   result_col9[8] <= result_col9[7];
   result_col9[9] <= result_col9[8];
   result_col9[10] <= result_col9[9];
   result_col9[11] <= result_col9[10];
   result_col9[12] <= result_col9[11];
   result_col9[13] <= result_col9[12];
   result_col9[14] <= result_col9[13];
   result_col9[15] <= result_col9[14];
   result_col9[16] <= result_col9[15];
   result_col9[17] <= result_col9[16];
   result_col9[18] <= result_col9[17];
   result_col9[19] <= result_col9[18];
   result_col9[20] <= result_col9[19];
   result_col9[21] <= result_col9[20];
   result_col9[22] <= result_col9[21];
   result_col9[23] <= result_col9[22];
   result_col9[24] <= result_col9[23];
   result_col9[25] <= result_col9[24];
   result_col9[26] <= result_col9[25];
   result_col9[27] <= result_col9[26];
   result_col9[28] <= result_col9[27];
   result_col9[29] <= result_col9[28];
   result_col9[30] <= result_col9[29];
   result_col9[31] <= result_col9[30];
   result_col9[32] <= result_col9[31];
   result_col9[33] <= result_col9[32];
   result_col9[34] <= result_col9[33];
   result_col9[35] <= result_col9[34];
   result_col9[36] <= result_col9[35];
   result_col9[37] <= result_col9[36];
   result_col9[38] <= result_col9[37];
   result_col9[39] <= result_col9[38];
   result_col9[40] <= result_col9[39];
   result_col9[41] <= result_col9[40];
   result_col9[42] <= result_col9[41];
   result_col9[43] <= result_col9[42];
   result_col9[44] <= result_col9[43];
   result_col9[45] <= result_col9[44];
   result_col9[46] <= result_col9[45];
   result_col9[47] <= result_col9[46];
   result_col9[48] <= result_col9[47];
   result_col9[49] <= result_col9[48];
   result_col9[50] <= result_col9[49];
   result_col9[51] <= result_col9[50];
   result_col9[52] <= result_col9[51];
   result_col9[53] <= result_col9[52];
   result_col9[54] <= result_col9[53];
   result_col9[55] <= result_col9[54];
   result_col9[56] <= result_col9[55];
   result_col9[57] <= result_col9[56];
   result_col9[58] <= result_col9[57];
   result_col9[59] <= result_col9[58];
   result_col9[60] <= result_col9[59];
   result_col9[61] <= result_col9[60];
   result_col9[62] <= result_col9[61];
   result_col9[63] <= result_col9[62];
   result_col9[64] <= result_col9[63];
   result_col9[65] <= result_col9[64];
   result_col9[66] <= result_col9[65];
   result_col9[67] <= result_col9[66];
   result_col9[68] <= result_col9[67];
   result_col9[69] <= result_col9[68];
   result_col9[70] <= result_col9[69];
   result_col9[71] <= result_col9[70];
   result_col9[72] <= result_col9[71];
   result_col9[73] <= result_col9[72];
   result_col9[74] <= result_col9[73];
   result_col9[75] <= result_col9[74];
   result_col9[76] <= result_col9[75];
   result_col9[77] <= result_col9[76];
   result_col9[78] <= result_col9[77];
   result_col9[79] <= result_col9[78];
   result_col9[80] <= result_col9[79];
   result_col9[81] <= result_col9[80];
   result_col9[82] <= result_col9[81];
   result_col9[83] <= result_col9[82];
   result_col9[84] <= result_col9[83];
   result_col9[85] <= result_col9[84];
   result_col9[86] <= result_col9[85];
   result_col9[87] <= result_col9[86];
   result_col9[88] <= result_col9[87];
   result_col9[89] <= result_col9[88];
   result_col9[90] <= result_col9[89];
   result_col9[91] <= result_col9[90];

   result_col10[1] <= data_out_5_10;
   result_col10[2] <= result_col10[1];
   result_col10[3] <= result_col10[2];
   result_col10[4] <= result_col10[3];
   result_col10[5] <= result_col10[4];
   result_col10[6] <= result_col10[5];
   result_col10[7] <= result_col10[6];
   result_col10[8] <= result_col10[7];
   result_col10[9] <= result_col10[8];
   result_col10[10] <= result_col10[9];
   result_col10[11] <= result_col10[10];
   result_col10[12] <= result_col10[11];
   result_col10[13] <= result_col10[12];
   result_col10[14] <= result_col10[13];
   result_col10[15] <= result_col10[14];
   result_col10[16] <= result_col10[15];
   result_col10[17] <= result_col10[16];
   result_col10[18] <= result_col10[17];
   result_col10[19] <= result_col10[18];
   result_col10[20] <= result_col10[19];
   result_col10[21] <= result_col10[20];
   result_col10[22] <= result_col10[21];
   result_col10[23] <= result_col10[22];
   result_col10[24] <= result_col10[23];
   result_col10[25] <= result_col10[24];
   result_col10[26] <= result_col10[25];
   result_col10[27] <= result_col10[26];
   result_col10[28] <= result_col10[27];
   result_col10[29] <= result_col10[28];
   result_col10[30] <= result_col10[29];
   result_col10[31] <= result_col10[30];
   result_col10[32] <= result_col10[31];
   result_col10[33] <= result_col10[32];
   result_col10[34] <= result_col10[33];
   result_col10[35] <= result_col10[34];
   result_col10[36] <= result_col10[35];
   result_col10[37] <= result_col10[36];
   result_col10[38] <= result_col10[37];
   result_col10[39] <= result_col10[38];
   result_col10[40] <= result_col10[39];
   result_col10[41] <= result_col10[40];
   result_col10[42] <= result_col10[41];
   result_col10[43] <= result_col10[42];
   result_col10[44] <= result_col10[43];
   result_col10[45] <= result_col10[44];
   result_col10[46] <= result_col10[45];
   result_col10[47] <= result_col10[46];
   result_col10[48] <= result_col10[47];
   result_col10[49] <= result_col10[48];
   result_col10[50] <= result_col10[49];
   result_col10[51] <= result_col10[50];
   result_col10[52] <= result_col10[51];
   result_col10[53] <= result_col10[52];
   result_col10[54] <= result_col10[53];
   result_col10[55] <= result_col10[54];
   result_col10[56] <= result_col10[55];
   result_col10[57] <= result_col10[56];
   result_col10[58] <= result_col10[57];
   result_col10[59] <= result_col10[58];
   result_col10[60] <= result_col10[59];
   result_col10[61] <= result_col10[60];
   result_col10[62] <= result_col10[61];
   result_col10[63] <= result_col10[62];
   result_col10[64] <= result_col10[63];
   result_col10[65] <= result_col10[64];
   result_col10[66] <= result_col10[65];
   result_col10[67] <= result_col10[66];
   result_col10[68] <= result_col10[67];
   result_col10[69] <= result_col10[68];
   result_col10[70] <= result_col10[69];
   result_col10[71] <= result_col10[70];
   result_col10[72] <= result_col10[71];
   result_col10[73] <= result_col10[72];
   result_col10[74] <= result_col10[73];
   result_col10[75] <= result_col10[74];
   result_col10[76] <= result_col10[75];
   result_col10[77] <= result_col10[76];
   result_col10[78] <= result_col10[77];
   result_col10[79] <= result_col10[78];
   result_col10[80] <= result_col10[79];
   result_col10[81] <= result_col10[80];
   result_col10[82] <= result_col10[81];
   result_col10[83] <= result_col10[82];
   result_col10[84] <= result_col10[83];
   result_col10[85] <= result_col10[84];
   result_col10[86] <= result_col10[85];
   result_col10[87] <= result_col10[86];
   result_col10[88] <= result_col10[87];
   result_col10[89] <= result_col10[88];
   result_col10[90] <= result_col10[89];

   result_col11[1] <= data_out_5_11;
   result_col11[2] <= result_col11[1];
   result_col11[3] <= result_col11[2];
   result_col11[4] <= result_col11[3];
   result_col11[5] <= result_col11[4];
   result_col11[6] <= result_col11[5];
   result_col11[7] <= result_col11[6];
   result_col11[8] <= result_col11[7];
   result_col11[9] <= result_col11[8];
   result_col11[10] <= result_col11[9];
   result_col11[11] <= result_col11[10];
   result_col11[12] <= result_col11[11];
   result_col11[13] <= result_col11[12];
   result_col11[14] <= result_col11[13];
   result_col11[15] <= result_col11[14];
   result_col11[16] <= result_col11[15];
   result_col11[17] <= result_col11[16];
   result_col11[18] <= result_col11[17];
   result_col11[19] <= result_col11[18];
   result_col11[20] <= result_col11[19];
   result_col11[21] <= result_col11[20];
   result_col11[22] <= result_col11[21];
   result_col11[23] <= result_col11[22];
   result_col11[24] <= result_col11[23];
   result_col11[25] <= result_col11[24];
   result_col11[26] <= result_col11[25];
   result_col11[27] <= result_col11[26];
   result_col11[28] <= result_col11[27];
   result_col11[29] <= result_col11[28];
   result_col11[30] <= result_col11[29];
   result_col11[31] <= result_col11[30];
   result_col11[32] <= result_col11[31];
   result_col11[33] <= result_col11[32];
   result_col11[34] <= result_col11[33];
   result_col11[35] <= result_col11[34];
   result_col11[36] <= result_col11[35];
   result_col11[37] <= result_col11[36];
   result_col11[38] <= result_col11[37];
   result_col11[39] <= result_col11[38];
   result_col11[40] <= result_col11[39];
   result_col11[41] <= result_col11[40];
   result_col11[42] <= result_col11[41];
   result_col11[43] <= result_col11[42];
   result_col11[44] <= result_col11[43];
   result_col11[45] <= result_col11[44];
   result_col11[46] <= result_col11[45];
   result_col11[47] <= result_col11[46];
   result_col11[48] <= result_col11[47];
   result_col11[49] <= result_col11[48];
   result_col11[50] <= result_col11[49];
   result_col11[51] <= result_col11[50];
   result_col11[52] <= result_col11[51];
   result_col11[53] <= result_col11[52];
   result_col11[54] <= result_col11[53];
   result_col11[55] <= result_col11[54];
   result_col11[56] <= result_col11[55];
   result_col11[57] <= result_col11[56];
   result_col11[58] <= result_col11[57];
   result_col11[59] <= result_col11[58];
   result_col11[60] <= result_col11[59];
   result_col11[61] <= result_col11[60];
   result_col11[62] <= result_col11[61];
   result_col11[63] <= result_col11[62];
   result_col11[64] <= result_col11[63];
   result_col11[65] <= result_col11[64];
   result_col11[66] <= result_col11[65];
   result_col11[67] <= result_col11[66];
   result_col11[68] <= result_col11[67];
   result_col11[69] <= result_col11[68];
   result_col11[70] <= result_col11[69];
   result_col11[71] <= result_col11[70];
   result_col11[72] <= result_col11[71];
   result_col11[73] <= result_col11[72];
   result_col11[74] <= result_col11[73];
   result_col11[75] <= result_col11[74];
   result_col11[76] <= result_col11[75];
   result_col11[77] <= result_col11[76];
   result_col11[78] <= result_col11[77];
   result_col11[79] <= result_col11[78];
   result_col11[80] <= result_col11[79];
   result_col11[81] <= result_col11[80];
   result_col11[82] <= result_col11[81];
   result_col11[83] <= result_col11[82];
   result_col11[84] <= result_col11[83];
   result_col11[85] <= result_col11[84];
   result_col11[86] <= result_col11[85];
   result_col11[87] <= result_col11[86];
   result_col11[88] <= result_col11[87];
   result_col11[89] <= result_col11[88];

   result_col12[1] <= data_out_5_12;
   result_col12[2] <= result_col12[1];
   result_col12[3] <= result_col12[2];
   result_col12[4] <= result_col12[3];
   result_col12[5] <= result_col12[4];
   result_col12[6] <= result_col12[5];
   result_col12[7] <= result_col12[6];
   result_col12[8] <= result_col12[7];
   result_col12[9] <= result_col12[8];
   result_col12[10] <= result_col12[9];
   result_col12[11] <= result_col12[10];
   result_col12[12] <= result_col12[11];
   result_col12[13] <= result_col12[12];
   result_col12[14] <= result_col12[13];
   result_col12[15] <= result_col12[14];
   result_col12[16] <= result_col12[15];
   result_col12[17] <= result_col12[16];
   result_col12[18] <= result_col12[17];
   result_col12[19] <= result_col12[18];
   result_col12[20] <= result_col12[19];
   result_col12[21] <= result_col12[20];
   result_col12[22] <= result_col12[21];
   result_col12[23] <= result_col12[22];
   result_col12[24] <= result_col12[23];
   result_col12[25] <= result_col12[24];
   result_col12[26] <= result_col12[25];
   result_col12[27] <= result_col12[26];
   result_col12[28] <= result_col12[27];
   result_col12[29] <= result_col12[28];
   result_col12[30] <= result_col12[29];
   result_col12[31] <= result_col12[30];
   result_col12[32] <= result_col12[31];
   result_col12[33] <= result_col12[32];
   result_col12[34] <= result_col12[33];
   result_col12[35] <= result_col12[34];
   result_col12[36] <= result_col12[35];
   result_col12[37] <= result_col12[36];
   result_col12[38] <= result_col12[37];
   result_col12[39] <= result_col12[38];
   result_col12[40] <= result_col12[39];
   result_col12[41] <= result_col12[40];
   result_col12[42] <= result_col12[41];
   result_col12[43] <= result_col12[42];
   result_col12[44] <= result_col12[43];
   result_col12[45] <= result_col12[44];
   result_col12[46] <= result_col12[45];
   result_col12[47] <= result_col12[46];
   result_col12[48] <= result_col12[47];
   result_col12[49] <= result_col12[48];
   result_col12[50] <= result_col12[49];
   result_col12[51] <= result_col12[50];
   result_col12[52] <= result_col12[51];
   result_col12[53] <= result_col12[52];
   result_col12[54] <= result_col12[53];
   result_col12[55] <= result_col12[54];
   result_col12[56] <= result_col12[55];
   result_col12[57] <= result_col12[56];
   result_col12[58] <= result_col12[57];
   result_col12[59] <= result_col12[58];
   result_col12[60] <= result_col12[59];
   result_col12[61] <= result_col12[60];
   result_col12[62] <= result_col12[61];
   result_col12[63] <= result_col12[62];
   result_col12[64] <= result_col12[63];
   result_col12[65] <= result_col12[64];
   result_col12[66] <= result_col12[65];
   result_col12[67] <= result_col12[66];
   result_col12[68] <= result_col12[67];
   result_col12[69] <= result_col12[68];
   result_col12[70] <= result_col12[69];
   result_col12[71] <= result_col12[70];
   result_col12[72] <= result_col12[71];
   result_col12[73] <= result_col12[72];
   result_col12[74] <= result_col12[73];
   result_col12[75] <= result_col12[74];
   result_col12[76] <= result_col12[75];
   result_col12[77] <= result_col12[76];
   result_col12[78] <= result_col12[77];
   result_col12[79] <= result_col12[78];
   result_col12[80] <= result_col12[79];
   result_col12[81] <= result_col12[80];
   result_col12[82] <= result_col12[81];
   result_col12[83] <= result_col12[82];
   result_col12[84] <= result_col12[83];
   result_col12[85] <= result_col12[84];
   result_col12[86] <= result_col12[85];
   result_col12[87] <= result_col12[86];
   result_col12[88] <= result_col12[87];

   result_col13[1] <= data_out_5_13;
   result_col13[2] <= result_col13[1];
   result_col13[3] <= result_col13[2];
   result_col13[4] <= result_col13[3];
   result_col13[5] <= result_col13[4];
   result_col13[6] <= result_col13[5];
   result_col13[7] <= result_col13[6];
   result_col13[8] <= result_col13[7];
   result_col13[9] <= result_col13[8];
   result_col13[10] <= result_col13[9];
   result_col13[11] <= result_col13[10];
   result_col13[12] <= result_col13[11];
   result_col13[13] <= result_col13[12];
   result_col13[14] <= result_col13[13];
   result_col13[15] <= result_col13[14];
   result_col13[16] <= result_col13[15];
   result_col13[17] <= result_col13[16];
   result_col13[18] <= result_col13[17];
   result_col13[19] <= result_col13[18];
   result_col13[20] <= result_col13[19];
   result_col13[21] <= result_col13[20];
   result_col13[22] <= result_col13[21];
   result_col13[23] <= result_col13[22];
   result_col13[24] <= result_col13[23];
   result_col13[25] <= result_col13[24];
   result_col13[26] <= result_col13[25];
   result_col13[27] <= result_col13[26];
   result_col13[28] <= result_col13[27];
   result_col13[29] <= result_col13[28];
   result_col13[30] <= result_col13[29];
   result_col13[31] <= result_col13[30];
   result_col13[32] <= result_col13[31];
   result_col13[33] <= result_col13[32];
   result_col13[34] <= result_col13[33];
   result_col13[35] <= result_col13[34];
   result_col13[36] <= result_col13[35];
   result_col13[37] <= result_col13[36];
   result_col13[38] <= result_col13[37];
   result_col13[39] <= result_col13[38];
   result_col13[40] <= result_col13[39];
   result_col13[41] <= result_col13[40];
   result_col13[42] <= result_col13[41];
   result_col13[43] <= result_col13[42];
   result_col13[44] <= result_col13[43];
   result_col13[45] <= result_col13[44];
   result_col13[46] <= result_col13[45];
   result_col13[47] <= result_col13[46];
   result_col13[48] <= result_col13[47];
   result_col13[49] <= result_col13[48];
   result_col13[50] <= result_col13[49];
   result_col13[51] <= result_col13[50];
   result_col13[52] <= result_col13[51];
   result_col13[53] <= result_col13[52];
   result_col13[54] <= result_col13[53];
   result_col13[55] <= result_col13[54];
   result_col13[56] <= result_col13[55];
   result_col13[57] <= result_col13[56];
   result_col13[58] <= result_col13[57];
   result_col13[59] <= result_col13[58];
   result_col13[60] <= result_col13[59];
   result_col13[61] <= result_col13[60];
   result_col13[62] <= result_col13[61];
   result_col13[63] <= result_col13[62];
   result_col13[64] <= result_col13[63];
   result_col13[65] <= result_col13[64];
   result_col13[66] <= result_col13[65];
   result_col13[67] <= result_col13[66];
   result_col13[68] <= result_col13[67];
   result_col13[69] <= result_col13[68];
   result_col13[70] <= result_col13[69];
   result_col13[71] <= result_col13[70];
   result_col13[72] <= result_col13[71];
   result_col13[73] <= result_col13[72];
   result_col13[74] <= result_col13[73];
   result_col13[75] <= result_col13[74];
   result_col13[76] <= result_col13[75];
   result_col13[77] <= result_col13[76];
   result_col13[78] <= result_col13[77];
   result_col13[79] <= result_col13[78];
   result_col13[80] <= result_col13[79];
   result_col13[81] <= result_col13[80];
   result_col13[82] <= result_col13[81];
   result_col13[83] <= result_col13[82];
   result_col13[84] <= result_col13[83];
   result_col13[85] <= result_col13[84];
   result_col13[86] <= result_col13[85];
   result_col13[87] <= result_col13[86];

   result_col14[1] <= data_out_5_14;
   result_col14[2] <= result_col14[1];
   result_col14[3] <= result_col14[2];
   result_col14[4] <= result_col14[3];
   result_col14[5] <= result_col14[4];
   result_col14[6] <= result_col14[5];
   result_col14[7] <= result_col14[6];
   result_col14[8] <= result_col14[7];
   result_col14[9] <= result_col14[8];
   result_col14[10] <= result_col14[9];
   result_col14[11] <= result_col14[10];
   result_col14[12] <= result_col14[11];
   result_col14[13] <= result_col14[12];
   result_col14[14] <= result_col14[13];
   result_col14[15] <= result_col14[14];
   result_col14[16] <= result_col14[15];
   result_col14[17] <= result_col14[16];
   result_col14[18] <= result_col14[17];
   result_col14[19] <= result_col14[18];
   result_col14[20] <= result_col14[19];
   result_col14[21] <= result_col14[20];
   result_col14[22] <= result_col14[21];
   result_col14[23] <= result_col14[22];
   result_col14[24] <= result_col14[23];
   result_col14[25] <= result_col14[24];
   result_col14[26] <= result_col14[25];
   result_col14[27] <= result_col14[26];
   result_col14[28] <= result_col14[27];
   result_col14[29] <= result_col14[28];
   result_col14[30] <= result_col14[29];
   result_col14[31] <= result_col14[30];
   result_col14[32] <= result_col14[31];
   result_col14[33] <= result_col14[32];
   result_col14[34] <= result_col14[33];
   result_col14[35] <= result_col14[34];
   result_col14[36] <= result_col14[35];
   result_col14[37] <= result_col14[36];
   result_col14[38] <= result_col14[37];
   result_col14[39] <= result_col14[38];
   result_col14[40] <= result_col14[39];
   result_col14[41] <= result_col14[40];
   result_col14[42] <= result_col14[41];
   result_col14[43] <= result_col14[42];
   result_col14[44] <= result_col14[43];
   result_col14[45] <= result_col14[44];
   result_col14[46] <= result_col14[45];
   result_col14[47] <= result_col14[46];
   result_col14[48] <= result_col14[47];
   result_col14[49] <= result_col14[48];
   result_col14[50] <= result_col14[49];
   result_col14[51] <= result_col14[50];
   result_col14[52] <= result_col14[51];
   result_col14[53] <= result_col14[52];
   result_col14[54] <= result_col14[53];
   result_col14[55] <= result_col14[54];
   result_col14[56] <= result_col14[55];
   result_col14[57] <= result_col14[56];
   result_col14[58] <= result_col14[57];
   result_col14[59] <= result_col14[58];
   result_col14[60] <= result_col14[59];
   result_col14[61] <= result_col14[60];
   result_col14[62] <= result_col14[61];
   result_col14[63] <= result_col14[62];
   result_col14[64] <= result_col14[63];
   result_col14[65] <= result_col14[64];
   result_col14[66] <= result_col14[65];
   result_col14[67] <= result_col14[66];
   result_col14[68] <= result_col14[67];
   result_col14[69] <= result_col14[68];
   result_col14[70] <= result_col14[69];
   result_col14[71] <= result_col14[70];
   result_col14[72] <= result_col14[71];
   result_col14[73] <= result_col14[72];
   result_col14[74] <= result_col14[73];
   result_col14[75] <= result_col14[74];
   result_col14[76] <= result_col14[75];
   result_col14[77] <= result_col14[76];
   result_col14[78] <= result_col14[77];
   result_col14[79] <= result_col14[78];
   result_col14[80] <= result_col14[79];
   result_col14[81] <= result_col14[80];
   result_col14[82] <= result_col14[81];
   result_col14[83] <= result_col14[82];
   result_col14[84] <= result_col14[83];
   result_col14[85] <= result_col14[84];
   result_col14[86] <= result_col14[85];

   result_col15[1] <= data_out_5_15;
   result_col15[2] <= result_col15[1];
   result_col15[3] <= result_col15[2];
   result_col15[4] <= result_col15[3];
   result_col15[5] <= result_col15[4];
   result_col15[6] <= result_col15[5];
   result_col15[7] <= result_col15[6];
   result_col15[8] <= result_col15[7];
   result_col15[9] <= result_col15[8];
   result_col15[10] <= result_col15[9];
   result_col15[11] <= result_col15[10];
   result_col15[12] <= result_col15[11];
   result_col15[13] <= result_col15[12];
   result_col15[14] <= result_col15[13];
   result_col15[15] <= result_col15[14];
   result_col15[16] <= result_col15[15];
   result_col15[17] <= result_col15[16];
   result_col15[18] <= result_col15[17];
   result_col15[19] <= result_col15[18];
   result_col15[20] <= result_col15[19];
   result_col15[21] <= result_col15[20];
   result_col15[22] <= result_col15[21];
   result_col15[23] <= result_col15[22];
   result_col15[24] <= result_col15[23];
   result_col15[25] <= result_col15[24];
   result_col15[26] <= result_col15[25];
   result_col15[27] <= result_col15[26];
   result_col15[28] <= result_col15[27];
   result_col15[29] <= result_col15[28];
   result_col15[30] <= result_col15[29];
   result_col15[31] <= result_col15[30];
   result_col15[32] <= result_col15[31];
   result_col15[33] <= result_col15[32];
   result_col15[34] <= result_col15[33];
   result_col15[35] <= result_col15[34];
   result_col15[36] <= result_col15[35];
   result_col15[37] <= result_col15[36];
   result_col15[38] <= result_col15[37];
   result_col15[39] <= result_col15[38];
   result_col15[40] <= result_col15[39];
   result_col15[41] <= result_col15[40];
   result_col15[42] <= result_col15[41];
   result_col15[43] <= result_col15[42];
   result_col15[44] <= result_col15[43];
   result_col15[45] <= result_col15[44];
   result_col15[46] <= result_col15[45];
   result_col15[47] <= result_col15[46];
   result_col15[48] <= result_col15[47];
   result_col15[49] <= result_col15[48];
   result_col15[50] <= result_col15[49];
   result_col15[51] <= result_col15[50];
   result_col15[52] <= result_col15[51];
   result_col15[53] <= result_col15[52];
   result_col15[54] <= result_col15[53];
   result_col15[55] <= result_col15[54];
   result_col15[56] <= result_col15[55];
   result_col15[57] <= result_col15[56];
   result_col15[58] <= result_col15[57];
   result_col15[59] <= result_col15[58];
   result_col15[60] <= result_col15[59];
   result_col15[61] <= result_col15[60];
   result_col15[62] <= result_col15[61];
   result_col15[63] <= result_col15[62];
   result_col15[64] <= result_col15[63];
   result_col15[65] <= result_col15[64];
   result_col15[66] <= result_col15[65];
   result_col15[67] <= result_col15[66];
   result_col15[68] <= result_col15[67];
   result_col15[69] <= result_col15[68];
   result_col15[70] <= result_col15[69];
   result_col15[71] <= result_col15[70];
   result_col15[72] <= result_col15[71];
   result_col15[73] <= result_col15[72];
   result_col15[74] <= result_col15[73];
   result_col15[75] <= result_col15[74];
   result_col15[76] <= result_col15[75];
   result_col15[77] <= result_col15[76];
   result_col15[78] <= result_col15[77];
   result_col15[79] <= result_col15[78];
   result_col15[80] <= result_col15[79];
   result_col15[81] <= result_col15[80];
   result_col15[82] <= result_col15[81];
   result_col15[83] <= result_col15[82];
   result_col15[84] <= result_col15[83];
   result_col15[85] <= result_col15[84];

   result_col16[1] <= data_out_5_16;
   result_col16[2] <= result_col16[1];
   result_col16[3] <= result_col16[2];
   result_col16[4] <= result_col16[3];
   result_col16[5] <= result_col16[4];
   result_col16[6] <= result_col16[5];
   result_col16[7] <= result_col16[6];
   result_col16[8] <= result_col16[7];
   result_col16[9] <= result_col16[8];
   result_col16[10] <= result_col16[9];
   result_col16[11] <= result_col16[10];
   result_col16[12] <= result_col16[11];
   result_col16[13] <= result_col16[12];
   result_col16[14] <= result_col16[13];
   result_col16[15] <= result_col16[14];
   result_col16[16] <= result_col16[15];
   result_col16[17] <= result_col16[16];
   result_col16[18] <= result_col16[17];
   result_col16[19] <= result_col16[18];
   result_col16[20] <= result_col16[19];
   result_col16[21] <= result_col16[20];
   result_col16[22] <= result_col16[21];
   result_col16[23] <= result_col16[22];
   result_col16[24] <= result_col16[23];
   result_col16[25] <= result_col16[24];
   result_col16[26] <= result_col16[25];
   result_col16[27] <= result_col16[26];
   result_col16[28] <= result_col16[27];
   result_col16[29] <= result_col16[28];
   result_col16[30] <= result_col16[29];
   result_col16[31] <= result_col16[30];
   result_col16[32] <= result_col16[31];
   result_col16[33] <= result_col16[32];
   result_col16[34] <= result_col16[33];
   result_col16[35] <= result_col16[34];
   result_col16[36] <= result_col16[35];
   result_col16[37] <= result_col16[36];
   result_col16[38] <= result_col16[37];
   result_col16[39] <= result_col16[38];
   result_col16[40] <= result_col16[39];
   result_col16[41] <= result_col16[40];
   result_col16[42] <= result_col16[41];
   result_col16[43] <= result_col16[42];
   result_col16[44] <= result_col16[43];
   result_col16[45] <= result_col16[44];
   result_col16[46] <= result_col16[45];
   result_col16[47] <= result_col16[46];
   result_col16[48] <= result_col16[47];
   result_col16[49] <= result_col16[48];
   result_col16[50] <= result_col16[49];
   result_col16[51] <= result_col16[50];
   result_col16[52] <= result_col16[51];
   result_col16[53] <= result_col16[52];
   result_col16[54] <= result_col16[53];
   result_col16[55] <= result_col16[54];
   result_col16[56] <= result_col16[55];
   result_col16[57] <= result_col16[56];
   result_col16[58] <= result_col16[57];
   result_col16[59] <= result_col16[58];
   result_col16[60] <= result_col16[59];
   result_col16[61] <= result_col16[60];
   result_col16[62] <= result_col16[61];
   result_col16[63] <= result_col16[62];
   result_col16[64] <= result_col16[63];
   result_col16[65] <= result_col16[64];
   result_col16[66] <= result_col16[65];
   result_col16[67] <= result_col16[66];
   result_col16[68] <= result_col16[67];
   result_col16[69] <= result_col16[68];
   result_col16[70] <= result_col16[69];
   result_col16[71] <= result_col16[70];
   result_col16[72] <= result_col16[71];
   result_col16[73] <= result_col16[72];
   result_col16[74] <= result_col16[73];
   result_col16[75] <= result_col16[74];
   result_col16[76] <= result_col16[75];
   result_col16[77] <= result_col16[76];
   result_col16[78] <= result_col16[77];
   result_col16[79] <= result_col16[78];
   result_col16[80] <= result_col16[79];
   result_col16[81] <= result_col16[80];
   result_col16[82] <= result_col16[81];
   result_col16[83] <= result_col16[82];
   result_col16[84] <= result_col16[83];

   result_col17[1] <= data_out_5_17;
   result_col17[2] <= result_col17[1];
   result_col17[3] <= result_col17[2];
   result_col17[4] <= result_col17[3];
   result_col17[5] <= result_col17[4];
   result_col17[6] <= result_col17[5];
   result_col17[7] <= result_col17[6];
   result_col17[8] <= result_col17[7];
   result_col17[9] <= result_col17[8];
   result_col17[10] <= result_col17[9];
   result_col17[11] <= result_col17[10];
   result_col17[12] <= result_col17[11];
   result_col17[13] <= result_col17[12];
   result_col17[14] <= result_col17[13];
   result_col17[15] <= result_col17[14];
   result_col17[16] <= result_col17[15];
   result_col17[17] <= result_col17[16];
   result_col17[18] <= result_col17[17];
   result_col17[19] <= result_col17[18];
   result_col17[20] <= result_col17[19];
   result_col17[21] <= result_col17[20];
   result_col17[22] <= result_col17[21];
   result_col17[23] <= result_col17[22];
   result_col17[24] <= result_col17[23];
   result_col17[25] <= result_col17[24];
   result_col17[26] <= result_col17[25];
   result_col17[27] <= result_col17[26];
   result_col17[28] <= result_col17[27];
   result_col17[29] <= result_col17[28];
   result_col17[30] <= result_col17[29];
   result_col17[31] <= result_col17[30];
   result_col17[32] <= result_col17[31];
   result_col17[33] <= result_col17[32];
   result_col17[34] <= result_col17[33];
   result_col17[35] <= result_col17[34];
   result_col17[36] <= result_col17[35];
   result_col17[37] <= result_col17[36];
   result_col17[38] <= result_col17[37];
   result_col17[39] <= result_col17[38];
   result_col17[40] <= result_col17[39];
   result_col17[41] <= result_col17[40];
   result_col17[42] <= result_col17[41];
   result_col17[43] <= result_col17[42];
   result_col17[44] <= result_col17[43];
   result_col17[45] <= result_col17[44];
   result_col17[46] <= result_col17[45];
   result_col17[47] <= result_col17[46];
   result_col17[48] <= result_col17[47];
   result_col17[49] <= result_col17[48];
   result_col17[50] <= result_col17[49];
   result_col17[51] <= result_col17[50];
   result_col17[52] <= result_col17[51];
   result_col17[53] <= result_col17[52];
   result_col17[54] <= result_col17[53];
   result_col17[55] <= result_col17[54];
   result_col17[56] <= result_col17[55];
   result_col17[57] <= result_col17[56];
   result_col17[58] <= result_col17[57];
   result_col17[59] <= result_col17[58];
   result_col17[60] <= result_col17[59];
   result_col17[61] <= result_col17[60];
   result_col17[62] <= result_col17[61];
   result_col17[63] <= result_col17[62];
   result_col17[64] <= result_col17[63];
   result_col17[65] <= result_col17[64];
   result_col17[66] <= result_col17[65];
   result_col17[67] <= result_col17[66];
   result_col17[68] <= result_col17[67];
   result_col17[69] <= result_col17[68];
   result_col17[70] <= result_col17[69];
   result_col17[71] <= result_col17[70];
   result_col17[72] <= result_col17[71];
   result_col17[73] <= result_col17[72];
   result_col17[74] <= result_col17[73];
   result_col17[75] <= result_col17[74];
   result_col17[76] <= result_col17[75];
   result_col17[77] <= result_col17[76];
   result_col17[78] <= result_col17[77];
   result_col17[79] <= result_col17[78];
   result_col17[80] <= result_col17[79];
   result_col17[81] <= result_col17[80];
   result_col17[82] <= result_col17[81];
   result_col17[83] <= result_col17[82];

   result_col18[1] <= data_out_5_18;
   result_col18[2] <= result_col18[1];
   result_col18[3] <= result_col18[2];
   result_col18[4] <= result_col18[3];
   result_col18[5] <= result_col18[4];
   result_col18[6] <= result_col18[5];
   result_col18[7] <= result_col18[6];
   result_col18[8] <= result_col18[7];
   result_col18[9] <= result_col18[8];
   result_col18[10] <= result_col18[9];
   result_col18[11] <= result_col18[10];
   result_col18[12] <= result_col18[11];
   result_col18[13] <= result_col18[12];
   result_col18[14] <= result_col18[13];
   result_col18[15] <= result_col18[14];
   result_col18[16] <= result_col18[15];
   result_col18[17] <= result_col18[16];
   result_col18[18] <= result_col18[17];
   result_col18[19] <= result_col18[18];
   result_col18[20] <= result_col18[19];
   result_col18[21] <= result_col18[20];
   result_col18[22] <= result_col18[21];
   result_col18[23] <= result_col18[22];
   result_col18[24] <= result_col18[23];
   result_col18[25] <= result_col18[24];
   result_col18[26] <= result_col18[25];
   result_col18[27] <= result_col18[26];
   result_col18[28] <= result_col18[27];
   result_col18[29] <= result_col18[28];
   result_col18[30] <= result_col18[29];
   result_col18[31] <= result_col18[30];
   result_col18[32] <= result_col18[31];
   result_col18[33] <= result_col18[32];
   result_col18[34] <= result_col18[33];
   result_col18[35] <= result_col18[34];
   result_col18[36] <= result_col18[35];
   result_col18[37] <= result_col18[36];
   result_col18[38] <= result_col18[37];
   result_col18[39] <= result_col18[38];
   result_col18[40] <= result_col18[39];
   result_col18[41] <= result_col18[40];
   result_col18[42] <= result_col18[41];
   result_col18[43] <= result_col18[42];
   result_col18[44] <= result_col18[43];
   result_col18[45] <= result_col18[44];
   result_col18[46] <= result_col18[45];
   result_col18[47] <= result_col18[46];
   result_col18[48] <= result_col18[47];
   result_col18[49] <= result_col18[48];
   result_col18[50] <= result_col18[49];
   result_col18[51] <= result_col18[50];
   result_col18[52] <= result_col18[51];
   result_col18[53] <= result_col18[52];
   result_col18[54] <= result_col18[53];
   result_col18[55] <= result_col18[54];
   result_col18[56] <= result_col18[55];
   result_col18[57] <= result_col18[56];
   result_col18[58] <= result_col18[57];
   result_col18[59] <= result_col18[58];
   result_col18[60] <= result_col18[59];
   result_col18[61] <= result_col18[60];
   result_col18[62] <= result_col18[61];
   result_col18[63] <= result_col18[62];
   result_col18[64] <= result_col18[63];
   result_col18[65] <= result_col18[64];
   result_col18[66] <= result_col18[65];
   result_col18[67] <= result_col18[66];
   result_col18[68] <= result_col18[67];
   result_col18[69] <= result_col18[68];
   result_col18[70] <= result_col18[69];
   result_col18[71] <= result_col18[70];
   result_col18[72] <= result_col18[71];
   result_col18[73] <= result_col18[72];
   result_col18[74] <= result_col18[73];
   result_col18[75] <= result_col18[74];
   result_col18[76] <= result_col18[75];
   result_col18[77] <= result_col18[76];
   result_col18[78] <= result_col18[77];
   result_col18[79] <= result_col18[78];
   result_col18[80] <= result_col18[79];
   result_col18[81] <= result_col18[80];
   result_col18[82] <= result_col18[81];

   result_col19[1] <= data_out_5_19;
   result_col19[2] <= result_col19[1];
   result_col19[3] <= result_col19[2];
   result_col19[4] <= result_col19[3];
   result_col19[5] <= result_col19[4];
   result_col19[6] <= result_col19[5];
   result_col19[7] <= result_col19[6];
   result_col19[8] <= result_col19[7];
   result_col19[9] <= result_col19[8];
   result_col19[10] <= result_col19[9];
   result_col19[11] <= result_col19[10];
   result_col19[12] <= result_col19[11];
   result_col19[13] <= result_col19[12];
   result_col19[14] <= result_col19[13];
   result_col19[15] <= result_col19[14];
   result_col19[16] <= result_col19[15];
   result_col19[17] <= result_col19[16];
   result_col19[18] <= result_col19[17];
   result_col19[19] <= result_col19[18];
   result_col19[20] <= result_col19[19];
   result_col19[21] <= result_col19[20];
   result_col19[22] <= result_col19[21];
   result_col19[23] <= result_col19[22];
   result_col19[24] <= result_col19[23];
   result_col19[25] <= result_col19[24];
   result_col19[26] <= result_col19[25];
   result_col19[27] <= result_col19[26];
   result_col19[28] <= result_col19[27];
   result_col19[29] <= result_col19[28];
   result_col19[30] <= result_col19[29];
   result_col19[31] <= result_col19[30];
   result_col19[32] <= result_col19[31];
   result_col19[33] <= result_col19[32];
   result_col19[34] <= result_col19[33];
   result_col19[35] <= result_col19[34];
   result_col19[36] <= result_col19[35];
   result_col19[37] <= result_col19[36];
   result_col19[38] <= result_col19[37];
   result_col19[39] <= result_col19[38];
   result_col19[40] <= result_col19[39];
   result_col19[41] <= result_col19[40];
   result_col19[42] <= result_col19[41];
   result_col19[43] <= result_col19[42];
   result_col19[44] <= result_col19[43];
   result_col19[45] <= result_col19[44];
   result_col19[46] <= result_col19[45];
   result_col19[47] <= result_col19[46];
   result_col19[48] <= result_col19[47];
   result_col19[49] <= result_col19[48];
   result_col19[50] <= result_col19[49];
   result_col19[51] <= result_col19[50];
   result_col19[52] <= result_col19[51];
   result_col19[53] <= result_col19[52];
   result_col19[54] <= result_col19[53];
   result_col19[55] <= result_col19[54];
   result_col19[56] <= result_col19[55];
   result_col19[57] <= result_col19[56];
   result_col19[58] <= result_col19[57];
   result_col19[59] <= result_col19[58];
   result_col19[60] <= result_col19[59];
   result_col19[61] <= result_col19[60];
   result_col19[62] <= result_col19[61];
   result_col19[63] <= result_col19[62];
   result_col19[64] <= result_col19[63];
   result_col19[65] <= result_col19[64];
   result_col19[66] <= result_col19[65];
   result_col19[67] <= result_col19[66];
   result_col19[68] <= result_col19[67];
   result_col19[69] <= result_col19[68];
   result_col19[70] <= result_col19[69];
   result_col19[71] <= result_col19[70];
   result_col19[72] <= result_col19[71];
   result_col19[73] <= result_col19[72];
   result_col19[74] <= result_col19[73];
   result_col19[75] <= result_col19[74];
   result_col19[76] <= result_col19[75];
   result_col19[77] <= result_col19[76];
   result_col19[78] <= result_col19[77];
   result_col19[79] <= result_col19[78];
   result_col19[80] <= result_col19[79];
   result_col19[81] <= result_col19[80];

   result_col20[1] <= data_out_5_20;
   result_col20[2] <= result_col20[1];
   result_col20[3] <= result_col20[2];
   result_col20[4] <= result_col20[3];
   result_col20[5] <= result_col20[4];
   result_col20[6] <= result_col20[5];
   result_col20[7] <= result_col20[6];
   result_col20[8] <= result_col20[7];
   result_col20[9] <= result_col20[8];
   result_col20[10] <= result_col20[9];
   result_col20[11] <= result_col20[10];
   result_col20[12] <= result_col20[11];
   result_col20[13] <= result_col20[12];
   result_col20[14] <= result_col20[13];
   result_col20[15] <= result_col20[14];
   result_col20[16] <= result_col20[15];
   result_col20[17] <= result_col20[16];
   result_col20[18] <= result_col20[17];
   result_col20[19] <= result_col20[18];
   result_col20[20] <= result_col20[19];
   result_col20[21] <= result_col20[20];
   result_col20[22] <= result_col20[21];
   result_col20[23] <= result_col20[22];
   result_col20[24] <= result_col20[23];
   result_col20[25] <= result_col20[24];
   result_col20[26] <= result_col20[25];
   result_col20[27] <= result_col20[26];
   result_col20[28] <= result_col20[27];
   result_col20[29] <= result_col20[28];
   result_col20[30] <= result_col20[29];
   result_col20[31] <= result_col20[30];
   result_col20[32] <= result_col20[31];
   result_col20[33] <= result_col20[32];
   result_col20[34] <= result_col20[33];
   result_col20[35] <= result_col20[34];
   result_col20[36] <= result_col20[35];
   result_col20[37] <= result_col20[36];
   result_col20[38] <= result_col20[37];
   result_col20[39] <= result_col20[38];
   result_col20[40] <= result_col20[39];
   result_col20[41] <= result_col20[40];
   result_col20[42] <= result_col20[41];
   result_col20[43] <= result_col20[42];
   result_col20[44] <= result_col20[43];
   result_col20[45] <= result_col20[44];
   result_col20[46] <= result_col20[45];
   result_col20[47] <= result_col20[46];
   result_col20[48] <= result_col20[47];
   result_col20[49] <= result_col20[48];
   result_col20[50] <= result_col20[49];
   result_col20[51] <= result_col20[50];
   result_col20[52] <= result_col20[51];
   result_col20[53] <= result_col20[52];
   result_col20[54] <= result_col20[53];
   result_col20[55] <= result_col20[54];
   result_col20[56] <= result_col20[55];
   result_col20[57] <= result_col20[56];
   result_col20[58] <= result_col20[57];
   result_col20[59] <= result_col20[58];
   result_col20[60] <= result_col20[59];
   result_col20[61] <= result_col20[60];
   result_col20[62] <= result_col20[61];
   result_col20[63] <= result_col20[62];
   result_col20[64] <= result_col20[63];
   result_col20[65] <= result_col20[64];
   result_col20[66] <= result_col20[65];
   result_col20[67] <= result_col20[66];
   result_col20[68] <= result_col20[67];
   result_col20[69] <= result_col20[68];
   result_col20[70] <= result_col20[69];
   result_col20[71] <= result_col20[70];
   result_col20[72] <= result_col20[71];
   result_col20[73] <= result_col20[72];
   result_col20[74] <= result_col20[73];
   result_col20[75] <= result_col20[74];
   result_col20[76] <= result_col20[75];
   result_col20[77] <= result_col20[76];
   result_col20[78] <= result_col20[77];
   result_col20[79] <= result_col20[78];
   result_col20[80] <= result_col20[79];

   result_col21[1] <= data_out_5_21;
   result_col21[2] <= result_col21[1];
   result_col21[3] <= result_col21[2];
   result_col21[4] <= result_col21[3];
   result_col21[5] <= result_col21[4];
   result_col21[6] <= result_col21[5];
   result_col21[7] <= result_col21[6];
   result_col21[8] <= result_col21[7];
   result_col21[9] <= result_col21[8];
   result_col21[10] <= result_col21[9];
   result_col21[11] <= result_col21[10];
   result_col21[12] <= result_col21[11];
   result_col21[13] <= result_col21[12];
   result_col21[14] <= result_col21[13];
   result_col21[15] <= result_col21[14];
   result_col21[16] <= result_col21[15];
   result_col21[17] <= result_col21[16];
   result_col21[18] <= result_col21[17];
   result_col21[19] <= result_col21[18];
   result_col21[20] <= result_col21[19];
   result_col21[21] <= result_col21[20];
   result_col21[22] <= result_col21[21];
   result_col21[23] <= result_col21[22];
   result_col21[24] <= result_col21[23];
   result_col21[25] <= result_col21[24];
   result_col21[26] <= result_col21[25];
   result_col21[27] <= result_col21[26];
   result_col21[28] <= result_col21[27];
   result_col21[29] <= result_col21[28];
   result_col21[30] <= result_col21[29];
   result_col21[31] <= result_col21[30];
   result_col21[32] <= result_col21[31];
   result_col21[33] <= result_col21[32];
   result_col21[34] <= result_col21[33];
   result_col21[35] <= result_col21[34];
   result_col21[36] <= result_col21[35];
   result_col21[37] <= result_col21[36];
   result_col21[38] <= result_col21[37];
   result_col21[39] <= result_col21[38];
   result_col21[40] <= result_col21[39];
   result_col21[41] <= result_col21[40];
   result_col21[42] <= result_col21[41];
   result_col21[43] <= result_col21[42];
   result_col21[44] <= result_col21[43];
   result_col21[45] <= result_col21[44];
   result_col21[46] <= result_col21[45];
   result_col21[47] <= result_col21[46];
   result_col21[48] <= result_col21[47];
   result_col21[49] <= result_col21[48];
   result_col21[50] <= result_col21[49];
   result_col21[51] <= result_col21[50];
   result_col21[52] <= result_col21[51];
   result_col21[53] <= result_col21[52];
   result_col21[54] <= result_col21[53];
   result_col21[55] <= result_col21[54];
   result_col21[56] <= result_col21[55];
   result_col21[57] <= result_col21[56];
   result_col21[58] <= result_col21[57];
   result_col21[59] <= result_col21[58];
   result_col21[60] <= result_col21[59];
   result_col21[61] <= result_col21[60];
   result_col21[62] <= result_col21[61];
   result_col21[63] <= result_col21[62];
   result_col21[64] <= result_col21[63];
   result_col21[65] <= result_col21[64];
   result_col21[66] <= result_col21[65];
   result_col21[67] <= result_col21[66];
   result_col21[68] <= result_col21[67];
   result_col21[69] <= result_col21[68];
   result_col21[70] <= result_col21[69];
   result_col21[71] <= result_col21[70];
   result_col21[72] <= result_col21[71];
   result_col21[73] <= result_col21[72];
   result_col21[74] <= result_col21[73];
   result_col21[75] <= result_col21[74];
   result_col21[76] <= result_col21[75];
   result_col21[77] <= result_col21[76];
   result_col21[78] <= result_col21[77];
   result_col21[79] <= result_col21[78];

   result_col22[1] <= data_out_5_22;
   result_col22[2] <= result_col22[1];
   result_col22[3] <= result_col22[2];
   result_col22[4] <= result_col22[3];
   result_col22[5] <= result_col22[4];
   result_col22[6] <= result_col22[5];
   result_col22[7] <= result_col22[6];
   result_col22[8] <= result_col22[7];
   result_col22[9] <= result_col22[8];
   result_col22[10] <= result_col22[9];
   result_col22[11] <= result_col22[10];
   result_col22[12] <= result_col22[11];
   result_col22[13] <= result_col22[12];
   result_col22[14] <= result_col22[13];
   result_col22[15] <= result_col22[14];
   result_col22[16] <= result_col22[15];
   result_col22[17] <= result_col22[16];
   result_col22[18] <= result_col22[17];
   result_col22[19] <= result_col22[18];
   result_col22[20] <= result_col22[19];
   result_col22[21] <= result_col22[20];
   result_col22[22] <= result_col22[21];
   result_col22[23] <= result_col22[22];
   result_col22[24] <= result_col22[23];
   result_col22[25] <= result_col22[24];
   result_col22[26] <= result_col22[25];
   result_col22[27] <= result_col22[26];
   result_col22[28] <= result_col22[27];
   result_col22[29] <= result_col22[28];
   result_col22[30] <= result_col22[29];
   result_col22[31] <= result_col22[30];
   result_col22[32] <= result_col22[31];
   result_col22[33] <= result_col22[32];
   result_col22[34] <= result_col22[33];
   result_col22[35] <= result_col22[34];
   result_col22[36] <= result_col22[35];
   result_col22[37] <= result_col22[36];
   result_col22[38] <= result_col22[37];
   result_col22[39] <= result_col22[38];
   result_col22[40] <= result_col22[39];
   result_col22[41] <= result_col22[40];
   result_col22[42] <= result_col22[41];
   result_col22[43] <= result_col22[42];
   result_col22[44] <= result_col22[43];
   result_col22[45] <= result_col22[44];
   result_col22[46] <= result_col22[45];
   result_col22[47] <= result_col22[46];
   result_col22[48] <= result_col22[47];
   result_col22[49] <= result_col22[48];
   result_col22[50] <= result_col22[49];
   result_col22[51] <= result_col22[50];
   result_col22[52] <= result_col22[51];
   result_col22[53] <= result_col22[52];
   result_col22[54] <= result_col22[53];
   result_col22[55] <= result_col22[54];
   result_col22[56] <= result_col22[55];
   result_col22[57] <= result_col22[56];
   result_col22[58] <= result_col22[57];
   result_col22[59] <= result_col22[58];
   result_col22[60] <= result_col22[59];
   result_col22[61] <= result_col22[60];
   result_col22[62] <= result_col22[61];
   result_col22[63] <= result_col22[62];
   result_col22[64] <= result_col22[63];
   result_col22[65] <= result_col22[64];
   result_col22[66] <= result_col22[65];
   result_col22[67] <= result_col22[66];
   result_col22[68] <= result_col22[67];
   result_col22[69] <= result_col22[68];
   result_col22[70] <= result_col22[69];
   result_col22[71] <= result_col22[70];
   result_col22[72] <= result_col22[71];
   result_col22[73] <= result_col22[72];
   result_col22[74] <= result_col22[73];
   result_col22[75] <= result_col22[74];
   result_col22[76] <= result_col22[75];
   result_col22[77] <= result_col22[76];
   result_col22[78] <= result_col22[77];

   result_col23[1] <= data_out_5_23;
   result_col23[2] <= result_col23[1];
   result_col23[3] <= result_col23[2];
   result_col23[4] <= result_col23[3];
   result_col23[5] <= result_col23[4];
   result_col23[6] <= result_col23[5];
   result_col23[7] <= result_col23[6];
   result_col23[8] <= result_col23[7];
   result_col23[9] <= result_col23[8];
   result_col23[10] <= result_col23[9];
   result_col23[11] <= result_col23[10];
   result_col23[12] <= result_col23[11];
   result_col23[13] <= result_col23[12];
   result_col23[14] <= result_col23[13];
   result_col23[15] <= result_col23[14];
   result_col23[16] <= result_col23[15];
   result_col23[17] <= result_col23[16];
   result_col23[18] <= result_col23[17];
   result_col23[19] <= result_col23[18];
   result_col23[20] <= result_col23[19];
   result_col23[21] <= result_col23[20];
   result_col23[22] <= result_col23[21];
   result_col23[23] <= result_col23[22];
   result_col23[24] <= result_col23[23];
   result_col23[25] <= result_col23[24];
   result_col23[26] <= result_col23[25];
   result_col23[27] <= result_col23[26];
   result_col23[28] <= result_col23[27];
   result_col23[29] <= result_col23[28];
   result_col23[30] <= result_col23[29];
   result_col23[31] <= result_col23[30];
   result_col23[32] <= result_col23[31];
   result_col23[33] <= result_col23[32];
   result_col23[34] <= result_col23[33];
   result_col23[35] <= result_col23[34];
   result_col23[36] <= result_col23[35];
   result_col23[37] <= result_col23[36];
   result_col23[38] <= result_col23[37];
   result_col23[39] <= result_col23[38];
   result_col23[40] <= result_col23[39];
   result_col23[41] <= result_col23[40];
   result_col23[42] <= result_col23[41];
   result_col23[43] <= result_col23[42];
   result_col23[44] <= result_col23[43];
   result_col23[45] <= result_col23[44];
   result_col23[46] <= result_col23[45];
   result_col23[47] <= result_col23[46];
   result_col23[48] <= result_col23[47];
   result_col23[49] <= result_col23[48];
   result_col23[50] <= result_col23[49];
   result_col23[51] <= result_col23[50];
   result_col23[52] <= result_col23[51];
   result_col23[53] <= result_col23[52];
   result_col23[54] <= result_col23[53];
   result_col23[55] <= result_col23[54];
   result_col23[56] <= result_col23[55];
   result_col23[57] <= result_col23[56];
   result_col23[58] <= result_col23[57];
   result_col23[59] <= result_col23[58];
   result_col23[60] <= result_col23[59];
   result_col23[61] <= result_col23[60];
   result_col23[62] <= result_col23[61];
   result_col23[63] <= result_col23[62];
   result_col23[64] <= result_col23[63];
   result_col23[65] <= result_col23[64];
   result_col23[66] <= result_col23[65];
   result_col23[67] <= result_col23[66];
   result_col23[68] <= result_col23[67];
   result_col23[69] <= result_col23[68];
   result_col23[70] <= result_col23[69];
   result_col23[71] <= result_col23[70];
   result_col23[72] <= result_col23[71];
   result_col23[73] <= result_col23[72];
   result_col23[74] <= result_col23[73];
   result_col23[75] <= result_col23[74];
   result_col23[76] <= result_col23[75];
   result_col23[77] <= result_col23[76];

   result_col24[1] <= data_out_5_24;
   result_col24[2] <= result_col24[1];
   result_col24[3] <= result_col24[2];
   result_col24[4] <= result_col24[3];
   result_col24[5] <= result_col24[4];
   result_col24[6] <= result_col24[5];
   result_col24[7] <= result_col24[6];
   result_col24[8] <= result_col24[7];
   result_col24[9] <= result_col24[8];
   result_col24[10] <= result_col24[9];
   result_col24[11] <= result_col24[10];
   result_col24[12] <= result_col24[11];
   result_col24[13] <= result_col24[12];
   result_col24[14] <= result_col24[13];
   result_col24[15] <= result_col24[14];
   result_col24[16] <= result_col24[15];
   result_col24[17] <= result_col24[16];
   result_col24[18] <= result_col24[17];
   result_col24[19] <= result_col24[18];
   result_col24[20] <= result_col24[19];
   result_col24[21] <= result_col24[20];
   result_col24[22] <= result_col24[21];
   result_col24[23] <= result_col24[22];
   result_col24[24] <= result_col24[23];
   result_col24[25] <= result_col24[24];
   result_col24[26] <= result_col24[25];
   result_col24[27] <= result_col24[26];
   result_col24[28] <= result_col24[27];
   result_col24[29] <= result_col24[28];
   result_col24[30] <= result_col24[29];
   result_col24[31] <= result_col24[30];
   result_col24[32] <= result_col24[31];
   result_col24[33] <= result_col24[32];
   result_col24[34] <= result_col24[33];
   result_col24[35] <= result_col24[34];
   result_col24[36] <= result_col24[35];
   result_col24[37] <= result_col24[36];
   result_col24[38] <= result_col24[37];
   result_col24[39] <= result_col24[38];
   result_col24[40] <= result_col24[39];
   result_col24[41] <= result_col24[40];
   result_col24[42] <= result_col24[41];
   result_col24[43] <= result_col24[42];
   result_col24[44] <= result_col24[43];
   result_col24[45] <= result_col24[44];
   result_col24[46] <= result_col24[45];
   result_col24[47] <= result_col24[46];
   result_col24[48] <= result_col24[47];
   result_col24[49] <= result_col24[48];
   result_col24[50] <= result_col24[49];
   result_col24[51] <= result_col24[50];
   result_col24[52] <= result_col24[51];
   result_col24[53] <= result_col24[52];
   result_col24[54] <= result_col24[53];
   result_col24[55] <= result_col24[54];
   result_col24[56] <= result_col24[55];
   result_col24[57] <= result_col24[56];
   result_col24[58] <= result_col24[57];
   result_col24[59] <= result_col24[58];
   result_col24[60] <= result_col24[59];
   result_col24[61] <= result_col24[60];
   result_col24[62] <= result_col24[61];
   result_col24[63] <= result_col24[62];
   result_col24[64] <= result_col24[63];
   result_col24[65] <= result_col24[64];
   result_col24[66] <= result_col24[65];
   result_col24[67] <= result_col24[66];
   result_col24[68] <= result_col24[67];
   result_col24[69] <= result_col24[68];
   result_col24[70] <= result_col24[69];
   result_col24[71] <= result_col24[70];
   result_col24[72] <= result_col24[71];
   result_col24[73] <= result_col24[72];
   result_col24[74] <= result_col24[73];
   result_col24[75] <= result_col24[74];
   result_col24[76] <= result_col24[75];

   result_col25[1] <= data_out_5_25;
   result_col25[2] <= result_col25[1];
   result_col25[3] <= result_col25[2];
   result_col25[4] <= result_col25[3];
   result_col25[5] <= result_col25[4];
   result_col25[6] <= result_col25[5];
   result_col25[7] <= result_col25[6];
   result_col25[8] <= result_col25[7];
   result_col25[9] <= result_col25[8];
   result_col25[10] <= result_col25[9];
   result_col25[11] <= result_col25[10];
   result_col25[12] <= result_col25[11];
   result_col25[13] <= result_col25[12];
   result_col25[14] <= result_col25[13];
   result_col25[15] <= result_col25[14];
   result_col25[16] <= result_col25[15];
   result_col25[17] <= result_col25[16];
   result_col25[18] <= result_col25[17];
   result_col25[19] <= result_col25[18];
   result_col25[20] <= result_col25[19];
   result_col25[21] <= result_col25[20];
   result_col25[22] <= result_col25[21];
   result_col25[23] <= result_col25[22];
   result_col25[24] <= result_col25[23];
   result_col25[25] <= result_col25[24];
   result_col25[26] <= result_col25[25];
   result_col25[27] <= result_col25[26];
   result_col25[28] <= result_col25[27];
   result_col25[29] <= result_col25[28];
   result_col25[30] <= result_col25[29];
   result_col25[31] <= result_col25[30];
   result_col25[32] <= result_col25[31];
   result_col25[33] <= result_col25[32];
   result_col25[34] <= result_col25[33];
   result_col25[35] <= result_col25[34];
   result_col25[36] <= result_col25[35];
   result_col25[37] <= result_col25[36];
   result_col25[38] <= result_col25[37];
   result_col25[39] <= result_col25[38];
   result_col25[40] <= result_col25[39];
   result_col25[41] <= result_col25[40];
   result_col25[42] <= result_col25[41];
   result_col25[43] <= result_col25[42];
   result_col25[44] <= result_col25[43];
   result_col25[45] <= result_col25[44];
   result_col25[46] <= result_col25[45];
   result_col25[47] <= result_col25[46];
   result_col25[48] <= result_col25[47];
   result_col25[49] <= result_col25[48];
   result_col25[50] <= result_col25[49];
   result_col25[51] <= result_col25[50];
   result_col25[52] <= result_col25[51];
   result_col25[53] <= result_col25[52];
   result_col25[54] <= result_col25[53];
   result_col25[55] <= result_col25[54];
   result_col25[56] <= result_col25[55];
   result_col25[57] <= result_col25[56];
   result_col25[58] <= result_col25[57];
   result_col25[59] <= result_col25[58];
   result_col25[60] <= result_col25[59];
   result_col25[61] <= result_col25[60];
   result_col25[62] <= result_col25[61];
   result_col25[63] <= result_col25[62];
   result_col25[64] <= result_col25[63];
   result_col25[65] <= result_col25[64];
   result_col25[66] <= result_col25[65];
   result_col25[67] <= result_col25[66];
   result_col25[68] <= result_col25[67];
   result_col25[69] <= result_col25[68];
   result_col25[70] <= result_col25[69];
   result_col25[71] <= result_col25[70];
   result_col25[72] <= result_col25[71];
   result_col25[73] <= result_col25[72];
   result_col25[74] <= result_col25[73];
   result_col25[75] <= result_col25[74];

   result_col26[1] <= data_out_5_26;
   result_col26[2] <= result_col26[1];
   result_col26[3] <= result_col26[2];
   result_col26[4] <= result_col26[3];
   result_col26[5] <= result_col26[4];
   result_col26[6] <= result_col26[5];
   result_col26[7] <= result_col26[6];
   result_col26[8] <= result_col26[7];
   result_col26[9] <= result_col26[8];
   result_col26[10] <= result_col26[9];
   result_col26[11] <= result_col26[10];
   result_col26[12] <= result_col26[11];
   result_col26[13] <= result_col26[12];
   result_col26[14] <= result_col26[13];
   result_col26[15] <= result_col26[14];
   result_col26[16] <= result_col26[15];
   result_col26[17] <= result_col26[16];
   result_col26[18] <= result_col26[17];
   result_col26[19] <= result_col26[18];
   result_col26[20] <= result_col26[19];
   result_col26[21] <= result_col26[20];
   result_col26[22] <= result_col26[21];
   result_col26[23] <= result_col26[22];
   result_col26[24] <= result_col26[23];
   result_col26[25] <= result_col26[24];
   result_col26[26] <= result_col26[25];
   result_col26[27] <= result_col26[26];
   result_col26[28] <= result_col26[27];
   result_col26[29] <= result_col26[28];
   result_col26[30] <= result_col26[29];
   result_col26[31] <= result_col26[30];
   result_col26[32] <= result_col26[31];
   result_col26[33] <= result_col26[32];
   result_col26[34] <= result_col26[33];
   result_col26[35] <= result_col26[34];
   result_col26[36] <= result_col26[35];
   result_col26[37] <= result_col26[36];
   result_col26[38] <= result_col26[37];
   result_col26[39] <= result_col26[38];
   result_col26[40] <= result_col26[39];
   result_col26[41] <= result_col26[40];
   result_col26[42] <= result_col26[41];
   result_col26[43] <= result_col26[42];
   result_col26[44] <= result_col26[43];
   result_col26[45] <= result_col26[44];
   result_col26[46] <= result_col26[45];
   result_col26[47] <= result_col26[46];
   result_col26[48] <= result_col26[47];
   result_col26[49] <= result_col26[48];
   result_col26[50] <= result_col26[49];
   result_col26[51] <= result_col26[50];
   result_col26[52] <= result_col26[51];
   result_col26[53] <= result_col26[52];
   result_col26[54] <= result_col26[53];
   result_col26[55] <= result_col26[54];
   result_col26[56] <= result_col26[55];
   result_col26[57] <= result_col26[56];
   result_col26[58] <= result_col26[57];
   result_col26[59] <= result_col26[58];
   result_col26[60] <= result_col26[59];
   result_col26[61] <= result_col26[60];
   result_col26[62] <= result_col26[61];
   result_col26[63] <= result_col26[62];
   result_col26[64] <= result_col26[63];
   result_col26[65] <= result_col26[64];
   result_col26[66] <= result_col26[65];
   result_col26[67] <= result_col26[66];
   result_col26[68] <= result_col26[67];
   result_col26[69] <= result_col26[68];
   result_col26[70] <= result_col26[69];
   result_col26[71] <= result_col26[70];
   result_col26[72] <= result_col26[71];
   result_col26[73] <= result_col26[72];
   result_col26[74] <= result_col26[73];

   result_col27[1] <= data_out_5_27;
   result_col27[2] <= result_col27[1];
   result_col27[3] <= result_col27[2];
   result_col27[4] <= result_col27[3];
   result_col27[5] <= result_col27[4];
   result_col27[6] <= result_col27[5];
   result_col27[7] <= result_col27[6];
   result_col27[8] <= result_col27[7];
   result_col27[9] <= result_col27[8];
   result_col27[10] <= result_col27[9];
   result_col27[11] <= result_col27[10];
   result_col27[12] <= result_col27[11];
   result_col27[13] <= result_col27[12];
   result_col27[14] <= result_col27[13];
   result_col27[15] <= result_col27[14];
   result_col27[16] <= result_col27[15];
   result_col27[17] <= result_col27[16];
   result_col27[18] <= result_col27[17];
   result_col27[19] <= result_col27[18];
   result_col27[20] <= result_col27[19];
   result_col27[21] <= result_col27[20];
   result_col27[22] <= result_col27[21];
   result_col27[23] <= result_col27[22];
   result_col27[24] <= result_col27[23];
   result_col27[25] <= result_col27[24];
   result_col27[26] <= result_col27[25];
   result_col27[27] <= result_col27[26];
   result_col27[28] <= result_col27[27];
   result_col27[29] <= result_col27[28];
   result_col27[30] <= result_col27[29];
   result_col27[31] <= result_col27[30];
   result_col27[32] <= result_col27[31];
   result_col27[33] <= result_col27[32];
   result_col27[34] <= result_col27[33];
   result_col27[35] <= result_col27[34];
   result_col27[36] <= result_col27[35];
   result_col27[37] <= result_col27[36];
   result_col27[38] <= result_col27[37];
   result_col27[39] <= result_col27[38];
   result_col27[40] <= result_col27[39];
   result_col27[41] <= result_col27[40];
   result_col27[42] <= result_col27[41];
   result_col27[43] <= result_col27[42];
   result_col27[44] <= result_col27[43];
   result_col27[45] <= result_col27[44];
   result_col27[46] <= result_col27[45];
   result_col27[47] <= result_col27[46];
   result_col27[48] <= result_col27[47];
   result_col27[49] <= result_col27[48];
   result_col27[50] <= result_col27[49];
   result_col27[51] <= result_col27[50];
   result_col27[52] <= result_col27[51];
   result_col27[53] <= result_col27[52];
   result_col27[54] <= result_col27[53];
   result_col27[55] <= result_col27[54];
   result_col27[56] <= result_col27[55];
   result_col27[57] <= result_col27[56];
   result_col27[58] <= result_col27[57];
   result_col27[59] <= result_col27[58];
   result_col27[60] <= result_col27[59];
   result_col27[61] <= result_col27[60];
   result_col27[62] <= result_col27[61];
   result_col27[63] <= result_col27[62];
   result_col27[64] <= result_col27[63];
   result_col27[65] <= result_col27[64];
   result_col27[66] <= result_col27[65];
   result_col27[67] <= result_col27[66];
   result_col27[68] <= result_col27[67];
   result_col27[69] <= result_col27[68];
   result_col27[70] <= result_col27[69];
   result_col27[71] <= result_col27[70];
   result_col27[72] <= result_col27[71];
   result_col27[73] <= result_col27[72];

   result_col28[1] <= data_out_5_28;
   result_col28[2] <= result_col28[1];
   result_col28[3] <= result_col28[2];
   result_col28[4] <= result_col28[3];
   result_col28[5] <= result_col28[4];
   result_col28[6] <= result_col28[5];
   result_col28[7] <= result_col28[6];
   result_col28[8] <= result_col28[7];
   result_col28[9] <= result_col28[8];
   result_col28[10] <= result_col28[9];
   result_col28[11] <= result_col28[10];
   result_col28[12] <= result_col28[11];
   result_col28[13] <= result_col28[12];
   result_col28[14] <= result_col28[13];
   result_col28[15] <= result_col28[14];
   result_col28[16] <= result_col28[15];
   result_col28[17] <= result_col28[16];
   result_col28[18] <= result_col28[17];
   result_col28[19] <= result_col28[18];
   result_col28[20] <= result_col28[19];
   result_col28[21] <= result_col28[20];
   result_col28[22] <= result_col28[21];
   result_col28[23] <= result_col28[22];
   result_col28[24] <= result_col28[23];
   result_col28[25] <= result_col28[24];
   result_col28[26] <= result_col28[25];
   result_col28[27] <= result_col28[26];
   result_col28[28] <= result_col28[27];
   result_col28[29] <= result_col28[28];
   result_col28[30] <= result_col28[29];
   result_col28[31] <= result_col28[30];
   result_col28[32] <= result_col28[31];
   result_col28[33] <= result_col28[32];
   result_col28[34] <= result_col28[33];
   result_col28[35] <= result_col28[34];
   result_col28[36] <= result_col28[35];
   result_col28[37] <= result_col28[36];
   result_col28[38] <= result_col28[37];
   result_col28[39] <= result_col28[38];
   result_col28[40] <= result_col28[39];
   result_col28[41] <= result_col28[40];
   result_col28[42] <= result_col28[41];
   result_col28[43] <= result_col28[42];
   result_col28[44] <= result_col28[43];
   result_col28[45] <= result_col28[44];
   result_col28[46] <= result_col28[45];
   result_col28[47] <= result_col28[46];
   result_col28[48] <= result_col28[47];
   result_col28[49] <= result_col28[48];
   result_col28[50] <= result_col28[49];
   result_col28[51] <= result_col28[50];
   result_col28[52] <= result_col28[51];
   result_col28[53] <= result_col28[52];
   result_col28[54] <= result_col28[53];
   result_col28[55] <= result_col28[54];
   result_col28[56] <= result_col28[55];
   result_col28[57] <= result_col28[56];
   result_col28[58] <= result_col28[57];
   result_col28[59] <= result_col28[58];
   result_col28[60] <= result_col28[59];
   result_col28[61] <= result_col28[60];
   result_col28[62] <= result_col28[61];
   result_col28[63] <= result_col28[62];
   result_col28[64] <= result_col28[63];
   result_col28[65] <= result_col28[64];
   result_col28[66] <= result_col28[65];
   result_col28[67] <= result_col28[66];
   result_col28[68] <= result_col28[67];
   result_col28[69] <= result_col28[68];
   result_col28[70] <= result_col28[69];
   result_col28[71] <= result_col28[70];
   result_col28[72] <= result_col28[71];

   result_col29[1] <= data_out_5_29;
   result_col29[2] <= result_col29[1];
   result_col29[3] <= result_col29[2];
   result_col29[4] <= result_col29[3];
   result_col29[5] <= result_col29[4];
   result_col29[6] <= result_col29[5];
   result_col29[7] <= result_col29[6];
   result_col29[8] <= result_col29[7];
   result_col29[9] <= result_col29[8];
   result_col29[10] <= result_col29[9];
   result_col29[11] <= result_col29[10];
   result_col29[12] <= result_col29[11];
   result_col29[13] <= result_col29[12];
   result_col29[14] <= result_col29[13];
   result_col29[15] <= result_col29[14];
   result_col29[16] <= result_col29[15];
   result_col29[17] <= result_col29[16];
   result_col29[18] <= result_col29[17];
   result_col29[19] <= result_col29[18];
   result_col29[20] <= result_col29[19];
   result_col29[21] <= result_col29[20];
   result_col29[22] <= result_col29[21];
   result_col29[23] <= result_col29[22];
   result_col29[24] <= result_col29[23];
   result_col29[25] <= result_col29[24];
   result_col29[26] <= result_col29[25];
   result_col29[27] <= result_col29[26];
   result_col29[28] <= result_col29[27];
   result_col29[29] <= result_col29[28];
   result_col29[30] <= result_col29[29];
   result_col29[31] <= result_col29[30];
   result_col29[32] <= result_col29[31];
   result_col29[33] <= result_col29[32];
   result_col29[34] <= result_col29[33];
   result_col29[35] <= result_col29[34];
   result_col29[36] <= result_col29[35];
   result_col29[37] <= result_col29[36];
   result_col29[38] <= result_col29[37];
   result_col29[39] <= result_col29[38];
   result_col29[40] <= result_col29[39];
   result_col29[41] <= result_col29[40];
   result_col29[42] <= result_col29[41];
   result_col29[43] <= result_col29[42];
   result_col29[44] <= result_col29[43];
   result_col29[45] <= result_col29[44];
   result_col29[46] <= result_col29[45];
   result_col29[47] <= result_col29[46];
   result_col29[48] <= result_col29[47];
   result_col29[49] <= result_col29[48];
   result_col29[50] <= result_col29[49];
   result_col29[51] <= result_col29[50];
   result_col29[52] <= result_col29[51];
   result_col29[53] <= result_col29[52];
   result_col29[54] <= result_col29[53];
   result_col29[55] <= result_col29[54];
   result_col29[56] <= result_col29[55];
   result_col29[57] <= result_col29[56];
   result_col29[58] <= result_col29[57];
   result_col29[59] <= result_col29[58];
   result_col29[60] <= result_col29[59];
   result_col29[61] <= result_col29[60];
   result_col29[62] <= result_col29[61];
   result_col29[63] <= result_col29[62];
   result_col29[64] <= result_col29[63];
   result_col29[65] <= result_col29[64];
   result_col29[66] <= result_col29[65];
   result_col29[67] <= result_col29[66];
   result_col29[68] <= result_col29[67];
   result_col29[69] <= result_col29[68];
   result_col29[70] <= result_col29[69];
   result_col29[71] <= result_col29[70];

   result_col30[1] <= data_out_5_30;
   result_col30[2] <= result_col30[1];
   result_col30[3] <= result_col30[2];
   result_col30[4] <= result_col30[3];
   result_col30[5] <= result_col30[4];
   result_col30[6] <= result_col30[5];
   result_col30[7] <= result_col30[6];
   result_col30[8] <= result_col30[7];
   result_col30[9] <= result_col30[8];
   result_col30[10] <= result_col30[9];
   result_col30[11] <= result_col30[10];
   result_col30[12] <= result_col30[11];
   result_col30[13] <= result_col30[12];
   result_col30[14] <= result_col30[13];
   result_col30[15] <= result_col30[14];
   result_col30[16] <= result_col30[15];
   result_col30[17] <= result_col30[16];
   result_col30[18] <= result_col30[17];
   result_col30[19] <= result_col30[18];
   result_col30[20] <= result_col30[19];
   result_col30[21] <= result_col30[20];
   result_col30[22] <= result_col30[21];
   result_col30[23] <= result_col30[22];
   result_col30[24] <= result_col30[23];
   result_col30[25] <= result_col30[24];
   result_col30[26] <= result_col30[25];
   result_col30[27] <= result_col30[26];
   result_col30[28] <= result_col30[27];
   result_col30[29] <= result_col30[28];
   result_col30[30] <= result_col30[29];
   result_col30[31] <= result_col30[30];
   result_col30[32] <= result_col30[31];
   result_col30[33] <= result_col30[32];
   result_col30[34] <= result_col30[33];
   result_col30[35] <= result_col30[34];
   result_col30[36] <= result_col30[35];
   result_col30[37] <= result_col30[36];
   result_col30[38] <= result_col30[37];
   result_col30[39] <= result_col30[38];
   result_col30[40] <= result_col30[39];
   result_col30[41] <= result_col30[40];
   result_col30[42] <= result_col30[41];
   result_col30[43] <= result_col30[42];
   result_col30[44] <= result_col30[43];
   result_col30[45] <= result_col30[44];
   result_col30[46] <= result_col30[45];
   result_col30[47] <= result_col30[46];
   result_col30[48] <= result_col30[47];
   result_col30[49] <= result_col30[48];
   result_col30[50] <= result_col30[49];
   result_col30[51] <= result_col30[50];
   result_col30[52] <= result_col30[51];
   result_col30[53] <= result_col30[52];
   result_col30[54] <= result_col30[53];
   result_col30[55] <= result_col30[54];
   result_col30[56] <= result_col30[55];
   result_col30[57] <= result_col30[56];
   result_col30[58] <= result_col30[57];
   result_col30[59] <= result_col30[58];
   result_col30[60] <= result_col30[59];
   result_col30[61] <= result_col30[60];
   result_col30[62] <= result_col30[61];
   result_col30[63] <= result_col30[62];
   result_col30[64] <= result_col30[63];
   result_col30[65] <= result_col30[64];
   result_col30[66] <= result_col30[65];
   result_col30[67] <= result_col30[66];
   result_col30[68] <= result_col30[67];
   result_col30[69] <= result_col30[68];
   result_col30[70] <= result_col30[69];

   result_col31[1] <= data_out_5_31;
   result_col31[2] <= result_col31[1];
   result_col31[3] <= result_col31[2];
   result_col31[4] <= result_col31[3];
   result_col31[5] <= result_col31[4];
   result_col31[6] <= result_col31[5];
   result_col31[7] <= result_col31[6];
   result_col31[8] <= result_col31[7];
   result_col31[9] <= result_col31[8];
   result_col31[10] <= result_col31[9];
   result_col31[11] <= result_col31[10];
   result_col31[12] <= result_col31[11];
   result_col31[13] <= result_col31[12];
   result_col31[14] <= result_col31[13];
   result_col31[15] <= result_col31[14];
   result_col31[16] <= result_col31[15];
   result_col31[17] <= result_col31[16];
   result_col31[18] <= result_col31[17];
   result_col31[19] <= result_col31[18];
   result_col31[20] <= result_col31[19];
   result_col31[21] <= result_col31[20];
   result_col31[22] <= result_col31[21];
   result_col31[23] <= result_col31[22];
   result_col31[24] <= result_col31[23];
   result_col31[25] <= result_col31[24];
   result_col31[26] <= result_col31[25];
   result_col31[27] <= result_col31[26];
   result_col31[28] <= result_col31[27];
   result_col31[29] <= result_col31[28];
   result_col31[30] <= result_col31[29];
   result_col31[31] <= result_col31[30];
   result_col31[32] <= result_col31[31];
   result_col31[33] <= result_col31[32];
   result_col31[34] <= result_col31[33];
   result_col31[35] <= result_col31[34];
   result_col31[36] <= result_col31[35];
   result_col31[37] <= result_col31[36];
   result_col31[38] <= result_col31[37];
   result_col31[39] <= result_col31[38];
   result_col31[40] <= result_col31[39];
   result_col31[41] <= result_col31[40];
   result_col31[42] <= result_col31[41];
   result_col31[43] <= result_col31[42];
   result_col31[44] <= result_col31[43];
   result_col31[45] <= result_col31[44];
   result_col31[46] <= result_col31[45];
   result_col31[47] <= result_col31[46];
   result_col31[48] <= result_col31[47];
   result_col31[49] <= result_col31[48];
   result_col31[50] <= result_col31[49];
   result_col31[51] <= result_col31[50];
   result_col31[52] <= result_col31[51];
   result_col31[53] <= result_col31[52];
   result_col31[54] <= result_col31[53];
   result_col31[55] <= result_col31[54];
   result_col31[56] <= result_col31[55];
   result_col31[57] <= result_col31[56];
   result_col31[58] <= result_col31[57];
   result_col31[59] <= result_col31[58];
   result_col31[60] <= result_col31[59];
   result_col31[61] <= result_col31[60];
   result_col31[62] <= result_col31[61];
   result_col31[63] <= result_col31[62];
   result_col31[64] <= result_col31[63];
   result_col31[65] <= result_col31[64];
   result_col31[66] <= result_col31[65];
   result_col31[67] <= result_col31[66];
   result_col31[68] <= result_col31[67];
   result_col31[69] <= result_col31[68];

   result_col32[1] <= data_out_5_32;
   result_col32[2] <= result_col32[1];
   result_col32[3] <= result_col32[2];
   result_col32[4] <= result_col32[3];
   result_col32[5] <= result_col32[4];
   result_col32[6] <= result_col32[5];
   result_col32[7] <= result_col32[6];
   result_col32[8] <= result_col32[7];
   result_col32[9] <= result_col32[8];
   result_col32[10] <= result_col32[9];
   result_col32[11] <= result_col32[10];
   result_col32[12] <= result_col32[11];
   result_col32[13] <= result_col32[12];
   result_col32[14] <= result_col32[13];
   result_col32[15] <= result_col32[14];
   result_col32[16] <= result_col32[15];
   result_col32[17] <= result_col32[16];
   result_col32[18] <= result_col32[17];
   result_col32[19] <= result_col32[18];
   result_col32[20] <= result_col32[19];
   result_col32[21] <= result_col32[20];
   result_col32[22] <= result_col32[21];
   result_col32[23] <= result_col32[22];
   result_col32[24] <= result_col32[23];
   result_col32[25] <= result_col32[24];
   result_col32[26] <= result_col32[25];
   result_col32[27] <= result_col32[26];
   result_col32[28] <= result_col32[27];
   result_col32[29] <= result_col32[28];
   result_col32[30] <= result_col32[29];
   result_col32[31] <= result_col32[30];
   result_col32[32] <= result_col32[31];
   result_col32[33] <= result_col32[32];
   result_col32[34] <= result_col32[33];
   result_col32[35] <= result_col32[34];
   result_col32[36] <= result_col32[35];
   result_col32[37] <= result_col32[36];
   result_col32[38] <= result_col32[37];
   result_col32[39] <= result_col32[38];
   result_col32[40] <= result_col32[39];
   result_col32[41] <= result_col32[40];
   result_col32[42] <= result_col32[41];
   result_col32[43] <= result_col32[42];
   result_col32[44] <= result_col32[43];
   result_col32[45] <= result_col32[44];
   result_col32[46] <= result_col32[45];
   result_col32[47] <= result_col32[46];
   result_col32[48] <= result_col32[47];
   result_col32[49] <= result_col32[48];
   result_col32[50] <= result_col32[49];
   result_col32[51] <= result_col32[50];
   result_col32[52] <= result_col32[51];
   result_col32[53] <= result_col32[52];
   result_col32[54] <= result_col32[53];
   result_col32[55] <= result_col32[54];
   result_col32[56] <= result_col32[55];
   result_col32[57] <= result_col32[56];
   result_col32[58] <= result_col32[57];
   result_col32[59] <= result_col32[58];
   result_col32[60] <= result_col32[59];
   result_col32[61] <= result_col32[60];
   result_col32[62] <= result_col32[61];
   result_col32[63] <= result_col32[62];
   result_col32[64] <= result_col32[63];
   result_col32[65] <= result_col32[64];
   result_col32[66] <= result_col32[65];
   result_col32[67] <= result_col32[66];
   result_col32[68] <= result_col32[67];

   result_col33[1] <= data_out_5_33;
   result_col33[2] <= result_col33[1];
   result_col33[3] <= result_col33[2];
   result_col33[4] <= result_col33[3];
   result_col33[5] <= result_col33[4];
   result_col33[6] <= result_col33[5];
   result_col33[7] <= result_col33[6];
   result_col33[8] <= result_col33[7];
   result_col33[9] <= result_col33[8];
   result_col33[10] <= result_col33[9];
   result_col33[11] <= result_col33[10];
   result_col33[12] <= result_col33[11];
   result_col33[13] <= result_col33[12];
   result_col33[14] <= result_col33[13];
   result_col33[15] <= result_col33[14];
   result_col33[16] <= result_col33[15];
   result_col33[17] <= result_col33[16];
   result_col33[18] <= result_col33[17];
   result_col33[19] <= result_col33[18];
   result_col33[20] <= result_col33[19];
   result_col33[21] <= result_col33[20];
   result_col33[22] <= result_col33[21];
   result_col33[23] <= result_col33[22];
   result_col33[24] <= result_col33[23];
   result_col33[25] <= result_col33[24];
   result_col33[26] <= result_col33[25];
   result_col33[27] <= result_col33[26];
   result_col33[28] <= result_col33[27];
   result_col33[29] <= result_col33[28];
   result_col33[30] <= result_col33[29];
   result_col33[31] <= result_col33[30];
   result_col33[32] <= result_col33[31];
   result_col33[33] <= result_col33[32];
   result_col33[34] <= result_col33[33];
   result_col33[35] <= result_col33[34];
   result_col33[36] <= result_col33[35];
   result_col33[37] <= result_col33[36];
   result_col33[38] <= result_col33[37];
   result_col33[39] <= result_col33[38];
   result_col33[40] <= result_col33[39];
   result_col33[41] <= result_col33[40];
   result_col33[42] <= result_col33[41];
   result_col33[43] <= result_col33[42];
   result_col33[44] <= result_col33[43];
   result_col33[45] <= result_col33[44];
   result_col33[46] <= result_col33[45];
   result_col33[47] <= result_col33[46];
   result_col33[48] <= result_col33[47];
   result_col33[49] <= result_col33[48];
   result_col33[50] <= result_col33[49];
   result_col33[51] <= result_col33[50];
   result_col33[52] <= result_col33[51];
   result_col33[53] <= result_col33[52];
   result_col33[54] <= result_col33[53];
   result_col33[55] <= result_col33[54];
   result_col33[56] <= result_col33[55];
   result_col33[57] <= result_col33[56];
   result_col33[58] <= result_col33[57];
   result_col33[59] <= result_col33[58];
   result_col33[60] <= result_col33[59];
   result_col33[61] <= result_col33[60];
   result_col33[62] <= result_col33[61];
   result_col33[63] <= result_col33[62];
   result_col33[64] <= result_col33[63];
   result_col33[65] <= result_col33[64];
   result_col33[66] <= result_col33[65];
   result_col33[67] <= result_col33[66];

   result_col34[1] <= data_out_5_34;
   result_col34[2] <= result_col34[1];
   result_col34[3] <= result_col34[2];
   result_col34[4] <= result_col34[3];
   result_col34[5] <= result_col34[4];
   result_col34[6] <= result_col34[5];
   result_col34[7] <= result_col34[6];
   result_col34[8] <= result_col34[7];
   result_col34[9] <= result_col34[8];
   result_col34[10] <= result_col34[9];
   result_col34[11] <= result_col34[10];
   result_col34[12] <= result_col34[11];
   result_col34[13] <= result_col34[12];
   result_col34[14] <= result_col34[13];
   result_col34[15] <= result_col34[14];
   result_col34[16] <= result_col34[15];
   result_col34[17] <= result_col34[16];
   result_col34[18] <= result_col34[17];
   result_col34[19] <= result_col34[18];
   result_col34[20] <= result_col34[19];
   result_col34[21] <= result_col34[20];
   result_col34[22] <= result_col34[21];
   result_col34[23] <= result_col34[22];
   result_col34[24] <= result_col34[23];
   result_col34[25] <= result_col34[24];
   result_col34[26] <= result_col34[25];
   result_col34[27] <= result_col34[26];
   result_col34[28] <= result_col34[27];
   result_col34[29] <= result_col34[28];
   result_col34[30] <= result_col34[29];
   result_col34[31] <= result_col34[30];
   result_col34[32] <= result_col34[31];
   result_col34[33] <= result_col34[32];
   result_col34[34] <= result_col34[33];
   result_col34[35] <= result_col34[34];
   result_col34[36] <= result_col34[35];
   result_col34[37] <= result_col34[36];
   result_col34[38] <= result_col34[37];
   result_col34[39] <= result_col34[38];
   result_col34[40] <= result_col34[39];
   result_col34[41] <= result_col34[40];
   result_col34[42] <= result_col34[41];
   result_col34[43] <= result_col34[42];
   result_col34[44] <= result_col34[43];
   result_col34[45] <= result_col34[44];
   result_col34[46] <= result_col34[45];
   result_col34[47] <= result_col34[46];
   result_col34[48] <= result_col34[47];
   result_col34[49] <= result_col34[48];
   result_col34[50] <= result_col34[49];
   result_col34[51] <= result_col34[50];
   result_col34[52] <= result_col34[51];
   result_col34[53] <= result_col34[52];
   result_col34[54] <= result_col34[53];
   result_col34[55] <= result_col34[54];
   result_col34[56] <= result_col34[55];
   result_col34[57] <= result_col34[56];
   result_col34[58] <= result_col34[57];
   result_col34[59] <= result_col34[58];
   result_col34[60] <= result_col34[59];
   result_col34[61] <= result_col34[60];
   result_col34[62] <= result_col34[61];
   result_col34[63] <= result_col34[62];
   result_col34[64] <= result_col34[63];
   result_col34[65] <= result_col34[64];
   result_col34[66] <= result_col34[65];

   result_col35[1] <= data_out_5_35;
   result_col35[2] <= result_col35[1];
   result_col35[3] <= result_col35[2];
   result_col35[4] <= result_col35[3];
   result_col35[5] <= result_col35[4];
   result_col35[6] <= result_col35[5];
   result_col35[7] <= result_col35[6];
   result_col35[8] <= result_col35[7];
   result_col35[9] <= result_col35[8];
   result_col35[10] <= result_col35[9];
   result_col35[11] <= result_col35[10];
   result_col35[12] <= result_col35[11];
   result_col35[13] <= result_col35[12];
   result_col35[14] <= result_col35[13];
   result_col35[15] <= result_col35[14];
   result_col35[16] <= result_col35[15];
   result_col35[17] <= result_col35[16];
   result_col35[18] <= result_col35[17];
   result_col35[19] <= result_col35[18];
   result_col35[20] <= result_col35[19];
   result_col35[21] <= result_col35[20];
   result_col35[22] <= result_col35[21];
   result_col35[23] <= result_col35[22];
   result_col35[24] <= result_col35[23];
   result_col35[25] <= result_col35[24];
   result_col35[26] <= result_col35[25];
   result_col35[27] <= result_col35[26];
   result_col35[28] <= result_col35[27];
   result_col35[29] <= result_col35[28];
   result_col35[30] <= result_col35[29];
   result_col35[31] <= result_col35[30];
   result_col35[32] <= result_col35[31];
   result_col35[33] <= result_col35[32];
   result_col35[34] <= result_col35[33];
   result_col35[35] <= result_col35[34];
   result_col35[36] <= result_col35[35];
   result_col35[37] <= result_col35[36];
   result_col35[38] <= result_col35[37];
   result_col35[39] <= result_col35[38];
   result_col35[40] <= result_col35[39];
   result_col35[41] <= result_col35[40];
   result_col35[42] <= result_col35[41];
   result_col35[43] <= result_col35[42];
   result_col35[44] <= result_col35[43];
   result_col35[45] <= result_col35[44];
   result_col35[46] <= result_col35[45];
   result_col35[47] <= result_col35[46];
   result_col35[48] <= result_col35[47];
   result_col35[49] <= result_col35[48];
   result_col35[50] <= result_col35[49];
   result_col35[51] <= result_col35[50];
   result_col35[52] <= result_col35[51];
   result_col35[53] <= result_col35[52];
   result_col35[54] <= result_col35[53];
   result_col35[55] <= result_col35[54];
   result_col35[56] <= result_col35[55];
   result_col35[57] <= result_col35[56];
   result_col35[58] <= result_col35[57];
   result_col35[59] <= result_col35[58];
   result_col35[60] <= result_col35[59];
   result_col35[61] <= result_col35[60];
   result_col35[62] <= result_col35[61];
   result_col35[63] <= result_col35[62];
   result_col35[64] <= result_col35[63];
   result_col35[65] <= result_col35[64];

   result_col36[1] <= data_out_5_36;
   result_col36[2] <= result_col36[1];
   result_col36[3] <= result_col36[2];
   result_col36[4] <= result_col36[3];
   result_col36[5] <= result_col36[4];
   result_col36[6] <= result_col36[5];
   result_col36[7] <= result_col36[6];
   result_col36[8] <= result_col36[7];
   result_col36[9] <= result_col36[8];
   result_col36[10] <= result_col36[9];
   result_col36[11] <= result_col36[10];
   result_col36[12] <= result_col36[11];
   result_col36[13] <= result_col36[12];
   result_col36[14] <= result_col36[13];
   result_col36[15] <= result_col36[14];
   result_col36[16] <= result_col36[15];
   result_col36[17] <= result_col36[16];
   result_col36[18] <= result_col36[17];
   result_col36[19] <= result_col36[18];
   result_col36[20] <= result_col36[19];
   result_col36[21] <= result_col36[20];
   result_col36[22] <= result_col36[21];
   result_col36[23] <= result_col36[22];
   result_col36[24] <= result_col36[23];
   result_col36[25] <= result_col36[24];
   result_col36[26] <= result_col36[25];
   result_col36[27] <= result_col36[26];
   result_col36[28] <= result_col36[27];
   result_col36[29] <= result_col36[28];
   result_col36[30] <= result_col36[29];
   result_col36[31] <= result_col36[30];
   result_col36[32] <= result_col36[31];
   result_col36[33] <= result_col36[32];
   result_col36[34] <= result_col36[33];
   result_col36[35] <= result_col36[34];
   result_col36[36] <= result_col36[35];
   result_col36[37] <= result_col36[36];
   result_col36[38] <= result_col36[37];
   result_col36[39] <= result_col36[38];
   result_col36[40] <= result_col36[39];
   result_col36[41] <= result_col36[40];
   result_col36[42] <= result_col36[41];
   result_col36[43] <= result_col36[42];
   result_col36[44] <= result_col36[43];
   result_col36[45] <= result_col36[44];
   result_col36[46] <= result_col36[45];
   result_col36[47] <= result_col36[46];
   result_col36[48] <= result_col36[47];
   result_col36[49] <= result_col36[48];
   result_col36[50] <= result_col36[49];
   result_col36[51] <= result_col36[50];
   result_col36[52] <= result_col36[51];
   result_col36[53] <= result_col36[52];
   result_col36[54] <= result_col36[53];
   result_col36[55] <= result_col36[54];
   result_col36[56] <= result_col36[55];
   result_col36[57] <= result_col36[56];
   result_col36[58] <= result_col36[57];
   result_col36[59] <= result_col36[58];
   result_col36[60] <= result_col36[59];
   result_col36[61] <= result_col36[60];
   result_col36[62] <= result_col36[61];
   result_col36[63] <= result_col36[62];
   result_col36[64] <= result_col36[63];

   result_col37[1] <= data_out_5_37;
   result_col37[2] <= result_col37[1];
   result_col37[3] <= result_col37[2];
   result_col37[4] <= result_col37[3];
   result_col37[5] <= result_col37[4];
   result_col37[6] <= result_col37[5];
   result_col37[7] <= result_col37[6];
   result_col37[8] <= result_col37[7];
   result_col37[9] <= result_col37[8];
   result_col37[10] <= result_col37[9];
   result_col37[11] <= result_col37[10];
   result_col37[12] <= result_col37[11];
   result_col37[13] <= result_col37[12];
   result_col37[14] <= result_col37[13];
   result_col37[15] <= result_col37[14];
   result_col37[16] <= result_col37[15];
   result_col37[17] <= result_col37[16];
   result_col37[18] <= result_col37[17];
   result_col37[19] <= result_col37[18];
   result_col37[20] <= result_col37[19];
   result_col37[21] <= result_col37[20];
   result_col37[22] <= result_col37[21];
   result_col37[23] <= result_col37[22];
   result_col37[24] <= result_col37[23];
   result_col37[25] <= result_col37[24];
   result_col37[26] <= result_col37[25];
   result_col37[27] <= result_col37[26];
   result_col37[28] <= result_col37[27];
   result_col37[29] <= result_col37[28];
   result_col37[30] <= result_col37[29];
   result_col37[31] <= result_col37[30];
   result_col37[32] <= result_col37[31];
   result_col37[33] <= result_col37[32];
   result_col37[34] <= result_col37[33];
   result_col37[35] <= result_col37[34];
   result_col37[36] <= result_col37[35];
   result_col37[37] <= result_col37[36];
   result_col37[38] <= result_col37[37];
   result_col37[39] <= result_col37[38];
   result_col37[40] <= result_col37[39];
   result_col37[41] <= result_col37[40];
   result_col37[42] <= result_col37[41];
   result_col37[43] <= result_col37[42];
   result_col37[44] <= result_col37[43];
   result_col37[45] <= result_col37[44];
   result_col37[46] <= result_col37[45];
   result_col37[47] <= result_col37[46];
   result_col37[48] <= result_col37[47];
   result_col37[49] <= result_col37[48];
   result_col37[50] <= result_col37[49];
   result_col37[51] <= result_col37[50];
   result_col37[52] <= result_col37[51];
   result_col37[53] <= result_col37[52];
   result_col37[54] <= result_col37[53];
   result_col37[55] <= result_col37[54];
   result_col37[56] <= result_col37[55];
   result_col37[57] <= result_col37[56];
   result_col37[58] <= result_col37[57];
   result_col37[59] <= result_col37[58];
   result_col37[60] <= result_col37[59];
   result_col37[61] <= result_col37[60];
   result_col37[62] <= result_col37[61];
   result_col37[63] <= result_col37[62];

   result_col38[1] <= data_out_5_38;
   result_col38[2] <= result_col38[1];
   result_col38[3] <= result_col38[2];
   result_col38[4] <= result_col38[3];
   result_col38[5] <= result_col38[4];
   result_col38[6] <= result_col38[5];
   result_col38[7] <= result_col38[6];
   result_col38[8] <= result_col38[7];
   result_col38[9] <= result_col38[8];
   result_col38[10] <= result_col38[9];
   result_col38[11] <= result_col38[10];
   result_col38[12] <= result_col38[11];
   result_col38[13] <= result_col38[12];
   result_col38[14] <= result_col38[13];
   result_col38[15] <= result_col38[14];
   result_col38[16] <= result_col38[15];
   result_col38[17] <= result_col38[16];
   result_col38[18] <= result_col38[17];
   result_col38[19] <= result_col38[18];
   result_col38[20] <= result_col38[19];
   result_col38[21] <= result_col38[20];
   result_col38[22] <= result_col38[21];
   result_col38[23] <= result_col38[22];
   result_col38[24] <= result_col38[23];
   result_col38[25] <= result_col38[24];
   result_col38[26] <= result_col38[25];
   result_col38[27] <= result_col38[26];
   result_col38[28] <= result_col38[27];
   result_col38[29] <= result_col38[28];
   result_col38[30] <= result_col38[29];
   result_col38[31] <= result_col38[30];
   result_col38[32] <= result_col38[31];
   result_col38[33] <= result_col38[32];
   result_col38[34] <= result_col38[33];
   result_col38[35] <= result_col38[34];
   result_col38[36] <= result_col38[35];
   result_col38[37] <= result_col38[36];
   result_col38[38] <= result_col38[37];
   result_col38[39] <= result_col38[38];
   result_col38[40] <= result_col38[39];
   result_col38[41] <= result_col38[40];
   result_col38[42] <= result_col38[41];
   result_col38[43] <= result_col38[42];
   result_col38[44] <= result_col38[43];
   result_col38[45] <= result_col38[44];
   result_col38[46] <= result_col38[45];
   result_col38[47] <= result_col38[46];
   result_col38[48] <= result_col38[47];
   result_col38[49] <= result_col38[48];
   result_col38[50] <= result_col38[49];
   result_col38[51] <= result_col38[50];
   result_col38[52] <= result_col38[51];
   result_col38[53] <= result_col38[52];
   result_col38[54] <= result_col38[53];
   result_col38[55] <= result_col38[54];
   result_col38[56] <= result_col38[55];
   result_col38[57] <= result_col38[56];
   result_col38[58] <= result_col38[57];
   result_col38[59] <= result_col38[58];
   result_col38[60] <= result_col38[59];
   result_col38[61] <= result_col38[60];
   result_col38[62] <= result_col38[61];

   result_col39[1] <= data_out_5_39;
   result_col39[2] <= result_col39[1];
   result_col39[3] <= result_col39[2];
   result_col39[4] <= result_col39[3];
   result_col39[5] <= result_col39[4];
   result_col39[6] <= result_col39[5];
   result_col39[7] <= result_col39[6];
   result_col39[8] <= result_col39[7];
   result_col39[9] <= result_col39[8];
   result_col39[10] <= result_col39[9];
   result_col39[11] <= result_col39[10];
   result_col39[12] <= result_col39[11];
   result_col39[13] <= result_col39[12];
   result_col39[14] <= result_col39[13];
   result_col39[15] <= result_col39[14];
   result_col39[16] <= result_col39[15];
   result_col39[17] <= result_col39[16];
   result_col39[18] <= result_col39[17];
   result_col39[19] <= result_col39[18];
   result_col39[20] <= result_col39[19];
   result_col39[21] <= result_col39[20];
   result_col39[22] <= result_col39[21];
   result_col39[23] <= result_col39[22];
   result_col39[24] <= result_col39[23];
   result_col39[25] <= result_col39[24];
   result_col39[26] <= result_col39[25];
   result_col39[27] <= result_col39[26];
   result_col39[28] <= result_col39[27];
   result_col39[29] <= result_col39[28];
   result_col39[30] <= result_col39[29];
   result_col39[31] <= result_col39[30];
   result_col39[32] <= result_col39[31];
   result_col39[33] <= result_col39[32];
   result_col39[34] <= result_col39[33];
   result_col39[35] <= result_col39[34];
   result_col39[36] <= result_col39[35];
   result_col39[37] <= result_col39[36];
   result_col39[38] <= result_col39[37];
   result_col39[39] <= result_col39[38];
   result_col39[40] <= result_col39[39];
   result_col39[41] <= result_col39[40];
   result_col39[42] <= result_col39[41];
   result_col39[43] <= result_col39[42];
   result_col39[44] <= result_col39[43];
   result_col39[45] <= result_col39[44];
   result_col39[46] <= result_col39[45];
   result_col39[47] <= result_col39[46];
   result_col39[48] <= result_col39[47];
   result_col39[49] <= result_col39[48];
   result_col39[50] <= result_col39[49];
   result_col39[51] <= result_col39[50];
   result_col39[52] <= result_col39[51];
   result_col39[53] <= result_col39[52];
   result_col39[54] <= result_col39[53];
   result_col39[55] <= result_col39[54];
   result_col39[56] <= result_col39[55];
   result_col39[57] <= result_col39[56];
   result_col39[58] <= result_col39[57];
   result_col39[59] <= result_col39[58];
   result_col39[60] <= result_col39[59];
   result_col39[61] <= result_col39[60];

   result_col40[1] <= data_out_5_40;
   result_col40[2] <= result_col40[1];
   result_col40[3] <= result_col40[2];
   result_col40[4] <= result_col40[3];
   result_col40[5] <= result_col40[4];
   result_col40[6] <= result_col40[5];
   result_col40[7] <= result_col40[6];
   result_col40[8] <= result_col40[7];
   result_col40[9] <= result_col40[8];
   result_col40[10] <= result_col40[9];
   result_col40[11] <= result_col40[10];
   result_col40[12] <= result_col40[11];
   result_col40[13] <= result_col40[12];
   result_col40[14] <= result_col40[13];
   result_col40[15] <= result_col40[14];
   result_col40[16] <= result_col40[15];
   result_col40[17] <= result_col40[16];
   result_col40[18] <= result_col40[17];
   result_col40[19] <= result_col40[18];
   result_col40[20] <= result_col40[19];
   result_col40[21] <= result_col40[20];
   result_col40[22] <= result_col40[21];
   result_col40[23] <= result_col40[22];
   result_col40[24] <= result_col40[23];
   result_col40[25] <= result_col40[24];
   result_col40[26] <= result_col40[25];
   result_col40[27] <= result_col40[26];
   result_col40[28] <= result_col40[27];
   result_col40[29] <= result_col40[28];
   result_col40[30] <= result_col40[29];
   result_col40[31] <= result_col40[30];
   result_col40[32] <= result_col40[31];
   result_col40[33] <= result_col40[32];
   result_col40[34] <= result_col40[33];
   result_col40[35] <= result_col40[34];
   result_col40[36] <= result_col40[35];
   result_col40[37] <= result_col40[36];
   result_col40[38] <= result_col40[37];
   result_col40[39] <= result_col40[38];
   result_col40[40] <= result_col40[39];
   result_col40[41] <= result_col40[40];
   result_col40[42] <= result_col40[41];
   result_col40[43] <= result_col40[42];
   result_col40[44] <= result_col40[43];
   result_col40[45] <= result_col40[44];
   result_col40[46] <= result_col40[45];
   result_col40[47] <= result_col40[46];
   result_col40[48] <= result_col40[47];
   result_col40[49] <= result_col40[48];
   result_col40[50] <= result_col40[49];
   result_col40[51] <= result_col40[50];
   result_col40[52] <= result_col40[51];
   result_col40[53] <= result_col40[52];
   result_col40[54] <= result_col40[53];
   result_col40[55] <= result_col40[54];
   result_col40[56] <= result_col40[55];
   result_col40[57] <= result_col40[56];
   result_col40[58] <= result_col40[57];
   result_col40[59] <= result_col40[58];
   result_col40[60] <= result_col40[59];

   result_col41[1] <= data_out_5_41;
   result_col41[2] <= result_col41[1];
   result_col41[3] <= result_col41[2];
   result_col41[4] <= result_col41[3];
   result_col41[5] <= result_col41[4];
   result_col41[6] <= result_col41[5];
   result_col41[7] <= result_col41[6];
   result_col41[8] <= result_col41[7];
   result_col41[9] <= result_col41[8];
   result_col41[10] <= result_col41[9];
   result_col41[11] <= result_col41[10];
   result_col41[12] <= result_col41[11];
   result_col41[13] <= result_col41[12];
   result_col41[14] <= result_col41[13];
   result_col41[15] <= result_col41[14];
   result_col41[16] <= result_col41[15];
   result_col41[17] <= result_col41[16];
   result_col41[18] <= result_col41[17];
   result_col41[19] <= result_col41[18];
   result_col41[20] <= result_col41[19];
   result_col41[21] <= result_col41[20];
   result_col41[22] <= result_col41[21];
   result_col41[23] <= result_col41[22];
   result_col41[24] <= result_col41[23];
   result_col41[25] <= result_col41[24];
   result_col41[26] <= result_col41[25];
   result_col41[27] <= result_col41[26];
   result_col41[28] <= result_col41[27];
   result_col41[29] <= result_col41[28];
   result_col41[30] <= result_col41[29];
   result_col41[31] <= result_col41[30];
   result_col41[32] <= result_col41[31];
   result_col41[33] <= result_col41[32];
   result_col41[34] <= result_col41[33];
   result_col41[35] <= result_col41[34];
   result_col41[36] <= result_col41[35];
   result_col41[37] <= result_col41[36];
   result_col41[38] <= result_col41[37];
   result_col41[39] <= result_col41[38];
   result_col41[40] <= result_col41[39];
   result_col41[41] <= result_col41[40];
   result_col41[42] <= result_col41[41];
   result_col41[43] <= result_col41[42];
   result_col41[44] <= result_col41[43];
   result_col41[45] <= result_col41[44];
   result_col41[46] <= result_col41[45];
   result_col41[47] <= result_col41[46];
   result_col41[48] <= result_col41[47];
   result_col41[49] <= result_col41[48];
   result_col41[50] <= result_col41[49];
   result_col41[51] <= result_col41[50];
   result_col41[52] <= result_col41[51];
   result_col41[53] <= result_col41[52];
   result_col41[54] <= result_col41[53];
   result_col41[55] <= result_col41[54];
   result_col41[56] <= result_col41[55];
   result_col41[57] <= result_col41[56];
   result_col41[58] <= result_col41[57];
   result_col41[59] <= result_col41[58];

   result_col42[1] <= data_out_5_42;
   result_col42[2] <= result_col42[1];
   result_col42[3] <= result_col42[2];
   result_col42[4] <= result_col42[3];
   result_col42[5] <= result_col42[4];
   result_col42[6] <= result_col42[5];
   result_col42[7] <= result_col42[6];
   result_col42[8] <= result_col42[7];
   result_col42[9] <= result_col42[8];
   result_col42[10] <= result_col42[9];
   result_col42[11] <= result_col42[10];
   result_col42[12] <= result_col42[11];
   result_col42[13] <= result_col42[12];
   result_col42[14] <= result_col42[13];
   result_col42[15] <= result_col42[14];
   result_col42[16] <= result_col42[15];
   result_col42[17] <= result_col42[16];
   result_col42[18] <= result_col42[17];
   result_col42[19] <= result_col42[18];
   result_col42[20] <= result_col42[19];
   result_col42[21] <= result_col42[20];
   result_col42[22] <= result_col42[21];
   result_col42[23] <= result_col42[22];
   result_col42[24] <= result_col42[23];
   result_col42[25] <= result_col42[24];
   result_col42[26] <= result_col42[25];
   result_col42[27] <= result_col42[26];
   result_col42[28] <= result_col42[27];
   result_col42[29] <= result_col42[28];
   result_col42[30] <= result_col42[29];
   result_col42[31] <= result_col42[30];
   result_col42[32] <= result_col42[31];
   result_col42[33] <= result_col42[32];
   result_col42[34] <= result_col42[33];
   result_col42[35] <= result_col42[34];
   result_col42[36] <= result_col42[35];
   result_col42[37] <= result_col42[36];
   result_col42[38] <= result_col42[37];
   result_col42[39] <= result_col42[38];
   result_col42[40] <= result_col42[39];
   result_col42[41] <= result_col42[40];
   result_col42[42] <= result_col42[41];
   result_col42[43] <= result_col42[42];
   result_col42[44] <= result_col42[43];
   result_col42[45] <= result_col42[44];
   result_col42[46] <= result_col42[45];
   result_col42[47] <= result_col42[46];
   result_col42[48] <= result_col42[47];
   result_col42[49] <= result_col42[48];
   result_col42[50] <= result_col42[49];
   result_col42[51] <= result_col42[50];
   result_col42[52] <= result_col42[51];
   result_col42[53] <= result_col42[52];
   result_col42[54] <= result_col42[53];
   result_col42[55] <= result_col42[54];
   result_col42[56] <= result_col42[55];
   result_col42[57] <= result_col42[56];
   result_col42[58] <= result_col42[57];

   result_col43[1] <= data_out_5_43;
   result_col43[2] <= result_col43[1];
   result_col43[3] <= result_col43[2];
   result_col43[4] <= result_col43[3];
   result_col43[5] <= result_col43[4];
   result_col43[6] <= result_col43[5];
   result_col43[7] <= result_col43[6];
   result_col43[8] <= result_col43[7];
   result_col43[9] <= result_col43[8];
   result_col43[10] <= result_col43[9];
   result_col43[11] <= result_col43[10];
   result_col43[12] <= result_col43[11];
   result_col43[13] <= result_col43[12];
   result_col43[14] <= result_col43[13];
   result_col43[15] <= result_col43[14];
   result_col43[16] <= result_col43[15];
   result_col43[17] <= result_col43[16];
   result_col43[18] <= result_col43[17];
   result_col43[19] <= result_col43[18];
   result_col43[20] <= result_col43[19];
   result_col43[21] <= result_col43[20];
   result_col43[22] <= result_col43[21];
   result_col43[23] <= result_col43[22];
   result_col43[24] <= result_col43[23];
   result_col43[25] <= result_col43[24];
   result_col43[26] <= result_col43[25];
   result_col43[27] <= result_col43[26];
   result_col43[28] <= result_col43[27];
   result_col43[29] <= result_col43[28];
   result_col43[30] <= result_col43[29];
   result_col43[31] <= result_col43[30];
   result_col43[32] <= result_col43[31];
   result_col43[33] <= result_col43[32];
   result_col43[34] <= result_col43[33];
   result_col43[35] <= result_col43[34];
   result_col43[36] <= result_col43[35];
   result_col43[37] <= result_col43[36];
   result_col43[38] <= result_col43[37];
   result_col43[39] <= result_col43[38];
   result_col43[40] <= result_col43[39];
   result_col43[41] <= result_col43[40];
   result_col43[42] <= result_col43[41];
   result_col43[43] <= result_col43[42];
   result_col43[44] <= result_col43[43];
   result_col43[45] <= result_col43[44];
   result_col43[46] <= result_col43[45];
   result_col43[47] <= result_col43[46];
   result_col43[48] <= result_col43[47];
   result_col43[49] <= result_col43[48];
   result_col43[50] <= result_col43[49];
   result_col43[51] <= result_col43[50];
   result_col43[52] <= result_col43[51];
   result_col43[53] <= result_col43[52];
   result_col43[54] <= result_col43[53];
   result_col43[55] <= result_col43[54];
   result_col43[56] <= result_col43[55];
   result_col43[57] <= result_col43[56];

   result_col44[1] <= data_out_5_44;
   result_col44[2] <= result_col44[1];
   result_col44[3] <= result_col44[2];
   result_col44[4] <= result_col44[3];
   result_col44[5] <= result_col44[4];
   result_col44[6] <= result_col44[5];
   result_col44[7] <= result_col44[6];
   result_col44[8] <= result_col44[7];
   result_col44[9] <= result_col44[8];
   result_col44[10] <= result_col44[9];
   result_col44[11] <= result_col44[10];
   result_col44[12] <= result_col44[11];
   result_col44[13] <= result_col44[12];
   result_col44[14] <= result_col44[13];
   result_col44[15] <= result_col44[14];
   result_col44[16] <= result_col44[15];
   result_col44[17] <= result_col44[16];
   result_col44[18] <= result_col44[17];
   result_col44[19] <= result_col44[18];
   result_col44[20] <= result_col44[19];
   result_col44[21] <= result_col44[20];
   result_col44[22] <= result_col44[21];
   result_col44[23] <= result_col44[22];
   result_col44[24] <= result_col44[23];
   result_col44[25] <= result_col44[24];
   result_col44[26] <= result_col44[25];
   result_col44[27] <= result_col44[26];
   result_col44[28] <= result_col44[27];
   result_col44[29] <= result_col44[28];
   result_col44[30] <= result_col44[29];
   result_col44[31] <= result_col44[30];
   result_col44[32] <= result_col44[31];
   result_col44[33] <= result_col44[32];
   result_col44[34] <= result_col44[33];
   result_col44[35] <= result_col44[34];
   result_col44[36] <= result_col44[35];
   result_col44[37] <= result_col44[36];
   result_col44[38] <= result_col44[37];
   result_col44[39] <= result_col44[38];
   result_col44[40] <= result_col44[39];
   result_col44[41] <= result_col44[40];
   result_col44[42] <= result_col44[41];
   result_col44[43] <= result_col44[42];
   result_col44[44] <= result_col44[43];
   result_col44[45] <= result_col44[44];
   result_col44[46] <= result_col44[45];
   result_col44[47] <= result_col44[46];
   result_col44[48] <= result_col44[47];
   result_col44[49] <= result_col44[48];
   result_col44[50] <= result_col44[49];
   result_col44[51] <= result_col44[50];
   result_col44[52] <= result_col44[51];
   result_col44[53] <= result_col44[52];
   result_col44[54] <= result_col44[53];
   result_col44[55] <= result_col44[54];
   result_col44[56] <= result_col44[55];

   result_col45[1] <= data_out_5_45;
   result_col45[2] <= result_col45[1];
   result_col45[3] <= result_col45[2];
   result_col45[4] <= result_col45[3];
   result_col45[5] <= result_col45[4];
   result_col45[6] <= result_col45[5];
   result_col45[7] <= result_col45[6];
   result_col45[8] <= result_col45[7];
   result_col45[9] <= result_col45[8];
   result_col45[10] <= result_col45[9];
   result_col45[11] <= result_col45[10];
   result_col45[12] <= result_col45[11];
   result_col45[13] <= result_col45[12];
   result_col45[14] <= result_col45[13];
   result_col45[15] <= result_col45[14];
   result_col45[16] <= result_col45[15];
   result_col45[17] <= result_col45[16];
   result_col45[18] <= result_col45[17];
   result_col45[19] <= result_col45[18];
   result_col45[20] <= result_col45[19];
   result_col45[21] <= result_col45[20];
   result_col45[22] <= result_col45[21];
   result_col45[23] <= result_col45[22];
   result_col45[24] <= result_col45[23];
   result_col45[25] <= result_col45[24];
   result_col45[26] <= result_col45[25];
   result_col45[27] <= result_col45[26];
   result_col45[28] <= result_col45[27];
   result_col45[29] <= result_col45[28];
   result_col45[30] <= result_col45[29];
   result_col45[31] <= result_col45[30];
   result_col45[32] <= result_col45[31];
   result_col45[33] <= result_col45[32];
   result_col45[34] <= result_col45[33];
   result_col45[35] <= result_col45[34];
   result_col45[36] <= result_col45[35];
   result_col45[37] <= result_col45[36];
   result_col45[38] <= result_col45[37];
   result_col45[39] <= result_col45[38];
   result_col45[40] <= result_col45[39];
   result_col45[41] <= result_col45[40];
   result_col45[42] <= result_col45[41];
   result_col45[43] <= result_col45[42];
   result_col45[44] <= result_col45[43];
   result_col45[45] <= result_col45[44];
   result_col45[46] <= result_col45[45];
   result_col45[47] <= result_col45[46];
   result_col45[48] <= result_col45[47];
   result_col45[49] <= result_col45[48];
   result_col45[50] <= result_col45[49];
   result_col45[51] <= result_col45[50];
   result_col45[52] <= result_col45[51];
   result_col45[53] <= result_col45[52];
   result_col45[54] <= result_col45[53];
   result_col45[55] <= result_col45[54];

   result_col46[1] <= data_out_5_46;
   result_col46[2] <= result_col46[1];
   result_col46[3] <= result_col46[2];
   result_col46[4] <= result_col46[3];
   result_col46[5] <= result_col46[4];
   result_col46[6] <= result_col46[5];
   result_col46[7] <= result_col46[6];
   result_col46[8] <= result_col46[7];
   result_col46[9] <= result_col46[8];
   result_col46[10] <= result_col46[9];
   result_col46[11] <= result_col46[10];
   result_col46[12] <= result_col46[11];
   result_col46[13] <= result_col46[12];
   result_col46[14] <= result_col46[13];
   result_col46[15] <= result_col46[14];
   result_col46[16] <= result_col46[15];
   result_col46[17] <= result_col46[16];
   result_col46[18] <= result_col46[17];
   result_col46[19] <= result_col46[18];
   result_col46[20] <= result_col46[19];
   result_col46[21] <= result_col46[20];
   result_col46[22] <= result_col46[21];
   result_col46[23] <= result_col46[22];
   result_col46[24] <= result_col46[23];
   result_col46[25] <= result_col46[24];
   result_col46[26] <= result_col46[25];
   result_col46[27] <= result_col46[26];
   result_col46[28] <= result_col46[27];
   result_col46[29] <= result_col46[28];
   result_col46[30] <= result_col46[29];
   result_col46[31] <= result_col46[30];
   result_col46[32] <= result_col46[31];
   result_col46[33] <= result_col46[32];
   result_col46[34] <= result_col46[33];
   result_col46[35] <= result_col46[34];
   result_col46[36] <= result_col46[35];
   result_col46[37] <= result_col46[36];
   result_col46[38] <= result_col46[37];
   result_col46[39] <= result_col46[38];
   result_col46[40] <= result_col46[39];
   result_col46[41] <= result_col46[40];
   result_col46[42] <= result_col46[41];
   result_col46[43] <= result_col46[42];
   result_col46[44] <= result_col46[43];
   result_col46[45] <= result_col46[44];
   result_col46[46] <= result_col46[45];
   result_col46[47] <= result_col46[46];
   result_col46[48] <= result_col46[47];
   result_col46[49] <= result_col46[48];
   result_col46[50] <= result_col46[49];
   result_col46[51] <= result_col46[50];
   result_col46[52] <= result_col46[51];
   result_col46[53] <= result_col46[52];
   result_col46[54] <= result_col46[53];

   result_col47[1] <= data_out_5_47;
   result_col47[2] <= result_col47[1];
   result_col47[3] <= result_col47[2];
   result_col47[4] <= result_col47[3];
   result_col47[5] <= result_col47[4];
   result_col47[6] <= result_col47[5];
   result_col47[7] <= result_col47[6];
   result_col47[8] <= result_col47[7];
   result_col47[9] <= result_col47[8];
   result_col47[10] <= result_col47[9];
   result_col47[11] <= result_col47[10];
   result_col47[12] <= result_col47[11];
   result_col47[13] <= result_col47[12];
   result_col47[14] <= result_col47[13];
   result_col47[15] <= result_col47[14];
   result_col47[16] <= result_col47[15];
   result_col47[17] <= result_col47[16];
   result_col47[18] <= result_col47[17];
   result_col47[19] <= result_col47[18];
   result_col47[20] <= result_col47[19];
   result_col47[21] <= result_col47[20];
   result_col47[22] <= result_col47[21];
   result_col47[23] <= result_col47[22];
   result_col47[24] <= result_col47[23];
   result_col47[25] <= result_col47[24];
   result_col47[26] <= result_col47[25];
   result_col47[27] <= result_col47[26];
   result_col47[28] <= result_col47[27];
   result_col47[29] <= result_col47[28];
   result_col47[30] <= result_col47[29];
   result_col47[31] <= result_col47[30];
   result_col47[32] <= result_col47[31];
   result_col47[33] <= result_col47[32];
   result_col47[34] <= result_col47[33];
   result_col47[35] <= result_col47[34];
   result_col47[36] <= result_col47[35];
   result_col47[37] <= result_col47[36];
   result_col47[38] <= result_col47[37];
   result_col47[39] <= result_col47[38];
   result_col47[40] <= result_col47[39];
   result_col47[41] <= result_col47[40];
   result_col47[42] <= result_col47[41];
   result_col47[43] <= result_col47[42];
   result_col47[44] <= result_col47[43];
   result_col47[45] <= result_col47[44];
   result_col47[46] <= result_col47[45];
   result_col47[47] <= result_col47[46];
   result_col47[48] <= result_col47[47];
   result_col47[49] <= result_col47[48];
   result_col47[50] <= result_col47[49];
   result_col47[51] <= result_col47[50];
   result_col47[52] <= result_col47[51];
   result_col47[53] <= result_col47[52];

   result_col48[1] <= data_out_5_48;
   result_col48[2] <= result_col48[1];
   result_col48[3] <= result_col48[2];
   result_col48[4] <= result_col48[3];
   result_col48[5] <= result_col48[4];
   result_col48[6] <= result_col48[5];
   result_col48[7] <= result_col48[6];
   result_col48[8] <= result_col48[7];
   result_col48[9] <= result_col48[8];
   result_col48[10] <= result_col48[9];
   result_col48[11] <= result_col48[10];
   result_col48[12] <= result_col48[11];
   result_col48[13] <= result_col48[12];
   result_col48[14] <= result_col48[13];
   result_col48[15] <= result_col48[14];
   result_col48[16] <= result_col48[15];
   result_col48[17] <= result_col48[16];
   result_col48[18] <= result_col48[17];
   result_col48[19] <= result_col48[18];
   result_col48[20] <= result_col48[19];
   result_col48[21] <= result_col48[20];
   result_col48[22] <= result_col48[21];
   result_col48[23] <= result_col48[22];
   result_col48[24] <= result_col48[23];
   result_col48[25] <= result_col48[24];
   result_col48[26] <= result_col48[25];
   result_col48[27] <= result_col48[26];
   result_col48[28] <= result_col48[27];
   result_col48[29] <= result_col48[28];
   result_col48[30] <= result_col48[29];
   result_col48[31] <= result_col48[30];
   result_col48[32] <= result_col48[31];
   result_col48[33] <= result_col48[32];
   result_col48[34] <= result_col48[33];
   result_col48[35] <= result_col48[34];
   result_col48[36] <= result_col48[35];
   result_col48[37] <= result_col48[36];
   result_col48[38] <= result_col48[37];
   result_col48[39] <= result_col48[38];
   result_col48[40] <= result_col48[39];
   result_col48[41] <= result_col48[40];
   result_col48[42] <= result_col48[41];
   result_col48[43] <= result_col48[42];
   result_col48[44] <= result_col48[43];
   result_col48[45] <= result_col48[44];
   result_col48[46] <= result_col48[45];
   result_col48[47] <= result_col48[46];
   result_col48[48] <= result_col48[47];
   result_col48[49] <= result_col48[48];
   result_col48[50] <= result_col48[49];
   result_col48[51] <= result_col48[50];
   result_col48[52] <= result_col48[51];

   result_col49[1] <= data_out_5_49;
   result_col49[2] <= result_col49[1];
   result_col49[3] <= result_col49[2];
   result_col49[4] <= result_col49[3];
   result_col49[5] <= result_col49[4];
   result_col49[6] <= result_col49[5];
   result_col49[7] <= result_col49[6];
   result_col49[8] <= result_col49[7];
   result_col49[9] <= result_col49[8];
   result_col49[10] <= result_col49[9];
   result_col49[11] <= result_col49[10];
   result_col49[12] <= result_col49[11];
   result_col49[13] <= result_col49[12];
   result_col49[14] <= result_col49[13];
   result_col49[15] <= result_col49[14];
   result_col49[16] <= result_col49[15];
   result_col49[17] <= result_col49[16];
   result_col49[18] <= result_col49[17];
   result_col49[19] <= result_col49[18];
   result_col49[20] <= result_col49[19];
   result_col49[21] <= result_col49[20];
   result_col49[22] <= result_col49[21];
   result_col49[23] <= result_col49[22];
   result_col49[24] <= result_col49[23];
   result_col49[25] <= result_col49[24];
   result_col49[26] <= result_col49[25];
   result_col49[27] <= result_col49[26];
   result_col49[28] <= result_col49[27];
   result_col49[29] <= result_col49[28];
   result_col49[30] <= result_col49[29];
   result_col49[31] <= result_col49[30];
   result_col49[32] <= result_col49[31];
   result_col49[33] <= result_col49[32];
   result_col49[34] <= result_col49[33];
   result_col49[35] <= result_col49[34];
   result_col49[36] <= result_col49[35];
   result_col49[37] <= result_col49[36];
   result_col49[38] <= result_col49[37];
   result_col49[39] <= result_col49[38];
   result_col49[40] <= result_col49[39];
   result_col49[41] <= result_col49[40];
   result_col49[42] <= result_col49[41];
   result_col49[43] <= result_col49[42];
   result_col49[44] <= result_col49[43];
   result_col49[45] <= result_col49[44];
   result_col49[46] <= result_col49[45];
   result_col49[47] <= result_col49[46];
   result_col49[48] <= result_col49[47];
   result_col49[49] <= result_col49[48];
   result_col49[50] <= result_col49[49];
   result_col49[51] <= result_col49[50];

   result_col50[1] <= data_out_5_50;
   result_col50[2] <= result_col50[1];
   result_col50[3] <= result_col50[2];
   result_col50[4] <= result_col50[3];
   result_col50[5] <= result_col50[4];
   result_col50[6] <= result_col50[5];
   result_col50[7] <= result_col50[6];
   result_col50[8] <= result_col50[7];
   result_col50[9] <= result_col50[8];
   result_col50[10] <= result_col50[9];
   result_col50[11] <= result_col50[10];
   result_col50[12] <= result_col50[11];
   result_col50[13] <= result_col50[12];
   result_col50[14] <= result_col50[13];
   result_col50[15] <= result_col50[14];
   result_col50[16] <= result_col50[15];
   result_col50[17] <= result_col50[16];
   result_col50[18] <= result_col50[17];
   result_col50[19] <= result_col50[18];
   result_col50[20] <= result_col50[19];
   result_col50[21] <= result_col50[20];
   result_col50[22] <= result_col50[21];
   result_col50[23] <= result_col50[22];
   result_col50[24] <= result_col50[23];
   result_col50[25] <= result_col50[24];
   result_col50[26] <= result_col50[25];
   result_col50[27] <= result_col50[26];
   result_col50[28] <= result_col50[27];
   result_col50[29] <= result_col50[28];
   result_col50[30] <= result_col50[29];
   result_col50[31] <= result_col50[30];
   result_col50[32] <= result_col50[31];
   result_col50[33] <= result_col50[32];
   result_col50[34] <= result_col50[33];
   result_col50[35] <= result_col50[34];
   result_col50[36] <= result_col50[35];
   result_col50[37] <= result_col50[36];
   result_col50[38] <= result_col50[37];
   result_col50[39] <= result_col50[38];
   result_col50[40] <= result_col50[39];
   result_col50[41] <= result_col50[40];
   result_col50[42] <= result_col50[41];
   result_col50[43] <= result_col50[42];
   result_col50[44] <= result_col50[43];
   result_col50[45] <= result_col50[44];
   result_col50[46] <= result_col50[45];
   result_col50[47] <= result_col50[46];
   result_col50[48] <= result_col50[47];
   result_col50[49] <= result_col50[48];
   result_col50[50] <= result_col50[49];

   result_col51[1] <= data_out_5_51;
   result_col51[2] <= result_col51[1];
   result_col51[3] <= result_col51[2];
   result_col51[4] <= result_col51[3];
   result_col51[5] <= result_col51[4];
   result_col51[6] <= result_col51[5];
   result_col51[7] <= result_col51[6];
   result_col51[8] <= result_col51[7];
   result_col51[9] <= result_col51[8];
   result_col51[10] <= result_col51[9];
   result_col51[11] <= result_col51[10];
   result_col51[12] <= result_col51[11];
   result_col51[13] <= result_col51[12];
   result_col51[14] <= result_col51[13];
   result_col51[15] <= result_col51[14];
   result_col51[16] <= result_col51[15];
   result_col51[17] <= result_col51[16];
   result_col51[18] <= result_col51[17];
   result_col51[19] <= result_col51[18];
   result_col51[20] <= result_col51[19];
   result_col51[21] <= result_col51[20];
   result_col51[22] <= result_col51[21];
   result_col51[23] <= result_col51[22];
   result_col51[24] <= result_col51[23];
   result_col51[25] <= result_col51[24];
   result_col51[26] <= result_col51[25];
   result_col51[27] <= result_col51[26];
   result_col51[28] <= result_col51[27];
   result_col51[29] <= result_col51[28];
   result_col51[30] <= result_col51[29];
   result_col51[31] <= result_col51[30];
   result_col51[32] <= result_col51[31];
   result_col51[33] <= result_col51[32];
   result_col51[34] <= result_col51[33];
   result_col51[35] <= result_col51[34];
   result_col51[36] <= result_col51[35];
   result_col51[37] <= result_col51[36];
   result_col51[38] <= result_col51[37];
   result_col51[39] <= result_col51[38];
   result_col51[40] <= result_col51[39];
   result_col51[41] <= result_col51[40];
   result_col51[42] <= result_col51[41];
   result_col51[43] <= result_col51[42];
   result_col51[44] <= result_col51[43];
   result_col51[45] <= result_col51[44];
   result_col51[46] <= result_col51[45];
   result_col51[47] <= result_col51[46];
   result_col51[48] <= result_col51[47];
   result_col51[49] <= result_col51[48];

   result_col52[1] <= data_out_5_52;
   result_col52[2] <= result_col52[1];
   result_col52[3] <= result_col52[2];
   result_col52[4] <= result_col52[3];
   result_col52[5] <= result_col52[4];
   result_col52[6] <= result_col52[5];
   result_col52[7] <= result_col52[6];
   result_col52[8] <= result_col52[7];
   result_col52[9] <= result_col52[8];
   result_col52[10] <= result_col52[9];
   result_col52[11] <= result_col52[10];
   result_col52[12] <= result_col52[11];
   result_col52[13] <= result_col52[12];
   result_col52[14] <= result_col52[13];
   result_col52[15] <= result_col52[14];
   result_col52[16] <= result_col52[15];
   result_col52[17] <= result_col52[16];
   result_col52[18] <= result_col52[17];
   result_col52[19] <= result_col52[18];
   result_col52[20] <= result_col52[19];
   result_col52[21] <= result_col52[20];
   result_col52[22] <= result_col52[21];
   result_col52[23] <= result_col52[22];
   result_col52[24] <= result_col52[23];
   result_col52[25] <= result_col52[24];
   result_col52[26] <= result_col52[25];
   result_col52[27] <= result_col52[26];
   result_col52[28] <= result_col52[27];
   result_col52[29] <= result_col52[28];
   result_col52[30] <= result_col52[29];
   result_col52[31] <= result_col52[30];
   result_col52[32] <= result_col52[31];
   result_col52[33] <= result_col52[32];
   result_col52[34] <= result_col52[33];
   result_col52[35] <= result_col52[34];
   result_col52[36] <= result_col52[35];
   result_col52[37] <= result_col52[36];
   result_col52[38] <= result_col52[37];
   result_col52[39] <= result_col52[38];
   result_col52[40] <= result_col52[39];
   result_col52[41] <= result_col52[40];
   result_col52[42] <= result_col52[41];
   result_col52[43] <= result_col52[42];
   result_col52[44] <= result_col52[43];
   result_col52[45] <= result_col52[44];
   result_col52[46] <= result_col52[45];
   result_col52[47] <= result_col52[46];
   result_col52[48] <= result_col52[47];

   result_col53[1] <= data_out_5_53;
   result_col53[2] <= result_col53[1];
   result_col53[3] <= result_col53[2];
   result_col53[4] <= result_col53[3];
   result_col53[5] <= result_col53[4];
   result_col53[6] <= result_col53[5];
   result_col53[7] <= result_col53[6];
   result_col53[8] <= result_col53[7];
   result_col53[9] <= result_col53[8];
   result_col53[10] <= result_col53[9];
   result_col53[11] <= result_col53[10];
   result_col53[12] <= result_col53[11];
   result_col53[13] <= result_col53[12];
   result_col53[14] <= result_col53[13];
   result_col53[15] <= result_col53[14];
   result_col53[16] <= result_col53[15];
   result_col53[17] <= result_col53[16];
   result_col53[18] <= result_col53[17];
   result_col53[19] <= result_col53[18];
   result_col53[20] <= result_col53[19];
   result_col53[21] <= result_col53[20];
   result_col53[22] <= result_col53[21];
   result_col53[23] <= result_col53[22];
   result_col53[24] <= result_col53[23];
   result_col53[25] <= result_col53[24];
   result_col53[26] <= result_col53[25];
   result_col53[27] <= result_col53[26];
   result_col53[28] <= result_col53[27];
   result_col53[29] <= result_col53[28];
   result_col53[30] <= result_col53[29];
   result_col53[31] <= result_col53[30];
   result_col53[32] <= result_col53[31];
   result_col53[33] <= result_col53[32];
   result_col53[34] <= result_col53[33];
   result_col53[35] <= result_col53[34];
   result_col53[36] <= result_col53[35];
   result_col53[37] <= result_col53[36];
   result_col53[38] <= result_col53[37];
   result_col53[39] <= result_col53[38];
   result_col53[40] <= result_col53[39];
   result_col53[41] <= result_col53[40];
   result_col53[42] <= result_col53[41];
   result_col53[43] <= result_col53[42];
   result_col53[44] <= result_col53[43];
   result_col53[45] <= result_col53[44];
   result_col53[46] <= result_col53[45];
   result_col53[47] <= result_col53[46];

   result_col54[1] <= data_out_5_54;
   result_col54[2] <= result_col54[1];
   result_col54[3] <= result_col54[2];
   result_col54[4] <= result_col54[3];
   result_col54[5] <= result_col54[4];
   result_col54[6] <= result_col54[5];
   result_col54[7] <= result_col54[6];
   result_col54[8] <= result_col54[7];
   result_col54[9] <= result_col54[8];
   result_col54[10] <= result_col54[9];
   result_col54[11] <= result_col54[10];
   result_col54[12] <= result_col54[11];
   result_col54[13] <= result_col54[12];
   result_col54[14] <= result_col54[13];
   result_col54[15] <= result_col54[14];
   result_col54[16] <= result_col54[15];
   result_col54[17] <= result_col54[16];
   result_col54[18] <= result_col54[17];
   result_col54[19] <= result_col54[18];
   result_col54[20] <= result_col54[19];
   result_col54[21] <= result_col54[20];
   result_col54[22] <= result_col54[21];
   result_col54[23] <= result_col54[22];
   result_col54[24] <= result_col54[23];
   result_col54[25] <= result_col54[24];
   result_col54[26] <= result_col54[25];
   result_col54[27] <= result_col54[26];
   result_col54[28] <= result_col54[27];
   result_col54[29] <= result_col54[28];
   result_col54[30] <= result_col54[29];
   result_col54[31] <= result_col54[30];
   result_col54[32] <= result_col54[31];
   result_col54[33] <= result_col54[32];
   result_col54[34] <= result_col54[33];
   result_col54[35] <= result_col54[34];
   result_col54[36] <= result_col54[35];
   result_col54[37] <= result_col54[36];
   result_col54[38] <= result_col54[37];
   result_col54[39] <= result_col54[38];
   result_col54[40] <= result_col54[39];
   result_col54[41] <= result_col54[40];
   result_col54[42] <= result_col54[41];
   result_col54[43] <= result_col54[42];
   result_col54[44] <= result_col54[43];
   result_col54[45] <= result_col54[44];
   result_col54[46] <= result_col54[45];

   result_col55[1] <= data_out_5_55;
   result_col55[2] <= result_col55[1];
   result_col55[3] <= result_col55[2];
   result_col55[4] <= result_col55[3];
   result_col55[5] <= result_col55[4];
   result_col55[6] <= result_col55[5];
   result_col55[7] <= result_col55[6];
   result_col55[8] <= result_col55[7];
   result_col55[9] <= result_col55[8];
   result_col55[10] <= result_col55[9];
   result_col55[11] <= result_col55[10];
   result_col55[12] <= result_col55[11];
   result_col55[13] <= result_col55[12];
   result_col55[14] <= result_col55[13];
   result_col55[15] <= result_col55[14];
   result_col55[16] <= result_col55[15];
   result_col55[17] <= result_col55[16];
   result_col55[18] <= result_col55[17];
   result_col55[19] <= result_col55[18];
   result_col55[20] <= result_col55[19];
   result_col55[21] <= result_col55[20];
   result_col55[22] <= result_col55[21];
   result_col55[23] <= result_col55[22];
   result_col55[24] <= result_col55[23];
   result_col55[25] <= result_col55[24];
   result_col55[26] <= result_col55[25];
   result_col55[27] <= result_col55[26];
   result_col55[28] <= result_col55[27];
   result_col55[29] <= result_col55[28];
   result_col55[30] <= result_col55[29];
   result_col55[31] <= result_col55[30];
   result_col55[32] <= result_col55[31];
   result_col55[33] <= result_col55[32];
   result_col55[34] <= result_col55[33];
   result_col55[35] <= result_col55[34];
   result_col55[36] <= result_col55[35];
   result_col55[37] <= result_col55[36];
   result_col55[38] <= result_col55[37];
   result_col55[39] <= result_col55[38];
   result_col55[40] <= result_col55[39];
   result_col55[41] <= result_col55[40];
   result_col55[42] <= result_col55[41];
   result_col55[43] <= result_col55[42];
   result_col55[44] <= result_col55[43];
   result_col55[45] <= result_col55[44];

   result_col56[1] <= data_out_5_56;
   result_col56[2] <= result_col56[1];
   result_col56[3] <= result_col56[2];
   result_col56[4] <= result_col56[3];
   result_col56[5] <= result_col56[4];
   result_col56[6] <= result_col56[5];
   result_col56[7] <= result_col56[6];
   result_col56[8] <= result_col56[7];
   result_col56[9] <= result_col56[8];
   result_col56[10] <= result_col56[9];
   result_col56[11] <= result_col56[10];
   result_col56[12] <= result_col56[11];
   result_col56[13] <= result_col56[12];
   result_col56[14] <= result_col56[13];
   result_col56[15] <= result_col56[14];
   result_col56[16] <= result_col56[15];
   result_col56[17] <= result_col56[16];
   result_col56[18] <= result_col56[17];
   result_col56[19] <= result_col56[18];
   result_col56[20] <= result_col56[19];
   result_col56[21] <= result_col56[20];
   result_col56[22] <= result_col56[21];
   result_col56[23] <= result_col56[22];
   result_col56[24] <= result_col56[23];
   result_col56[25] <= result_col56[24];
   result_col56[26] <= result_col56[25];
   result_col56[27] <= result_col56[26];
   result_col56[28] <= result_col56[27];
   result_col56[29] <= result_col56[28];
   result_col56[30] <= result_col56[29];
   result_col56[31] <= result_col56[30];
   result_col56[32] <= result_col56[31];
   result_col56[33] <= result_col56[32];
   result_col56[34] <= result_col56[33];
   result_col56[35] <= result_col56[34];
   result_col56[36] <= result_col56[35];
   result_col56[37] <= result_col56[36];
   result_col56[38] <= result_col56[37];
   result_col56[39] <= result_col56[38];
   result_col56[40] <= result_col56[39];
   result_col56[41] <= result_col56[40];
   result_col56[42] <= result_col56[41];
   result_col56[43] <= result_col56[42];
   result_col56[44] <= result_col56[43];

   result_col57[1] <= data_out_5_57;
   result_col57[2] <= result_col57[1];
   result_col57[3] <= result_col57[2];
   result_col57[4] <= result_col57[3];
   result_col57[5] <= result_col57[4];
   result_col57[6] <= result_col57[5];
   result_col57[7] <= result_col57[6];
   result_col57[8] <= result_col57[7];
   result_col57[9] <= result_col57[8];
   result_col57[10] <= result_col57[9];
   result_col57[11] <= result_col57[10];
   result_col57[12] <= result_col57[11];
   result_col57[13] <= result_col57[12];
   result_col57[14] <= result_col57[13];
   result_col57[15] <= result_col57[14];
   result_col57[16] <= result_col57[15];
   result_col57[17] <= result_col57[16];
   result_col57[18] <= result_col57[17];
   result_col57[19] <= result_col57[18];
   result_col57[20] <= result_col57[19];
   result_col57[21] <= result_col57[20];
   result_col57[22] <= result_col57[21];
   result_col57[23] <= result_col57[22];
   result_col57[24] <= result_col57[23];
   result_col57[25] <= result_col57[24];
   result_col57[26] <= result_col57[25];
   result_col57[27] <= result_col57[26];
   result_col57[28] <= result_col57[27];
   result_col57[29] <= result_col57[28];
   result_col57[30] <= result_col57[29];
   result_col57[31] <= result_col57[30];
   result_col57[32] <= result_col57[31];
   result_col57[33] <= result_col57[32];
   result_col57[34] <= result_col57[33];
   result_col57[35] <= result_col57[34];
   result_col57[36] <= result_col57[35];
   result_col57[37] <= result_col57[36];
   result_col57[38] <= result_col57[37];
   result_col57[39] <= result_col57[38];
   result_col57[40] <= result_col57[39];
   result_col57[41] <= result_col57[40];
   result_col57[42] <= result_col57[41];
   result_col57[43] <= result_col57[42];

   result_col58[1] <= data_out_5_58;
   result_col58[2] <= result_col58[1];
   result_col58[3] <= result_col58[2];
   result_col58[4] <= result_col58[3];
   result_col58[5] <= result_col58[4];
   result_col58[6] <= result_col58[5];
   result_col58[7] <= result_col58[6];
   result_col58[8] <= result_col58[7];
   result_col58[9] <= result_col58[8];
   result_col58[10] <= result_col58[9];
   result_col58[11] <= result_col58[10];
   result_col58[12] <= result_col58[11];
   result_col58[13] <= result_col58[12];
   result_col58[14] <= result_col58[13];
   result_col58[15] <= result_col58[14];
   result_col58[16] <= result_col58[15];
   result_col58[17] <= result_col58[16];
   result_col58[18] <= result_col58[17];
   result_col58[19] <= result_col58[18];
   result_col58[20] <= result_col58[19];
   result_col58[21] <= result_col58[20];
   result_col58[22] <= result_col58[21];
   result_col58[23] <= result_col58[22];
   result_col58[24] <= result_col58[23];
   result_col58[25] <= result_col58[24];
   result_col58[26] <= result_col58[25];
   result_col58[27] <= result_col58[26];
   result_col58[28] <= result_col58[27];
   result_col58[29] <= result_col58[28];
   result_col58[30] <= result_col58[29];
   result_col58[31] <= result_col58[30];
   result_col58[32] <= result_col58[31];
   result_col58[33] <= result_col58[32];
   result_col58[34] <= result_col58[33];
   result_col58[35] <= result_col58[34];
   result_col58[36] <= result_col58[35];
   result_col58[37] <= result_col58[36];
   result_col58[38] <= result_col58[37];
   result_col58[39] <= result_col58[38];
   result_col58[40] <= result_col58[39];
   result_col58[41] <= result_col58[40];
   result_col58[42] <= result_col58[41];

   result_col59[1] <= data_out_5_59;
   result_col59[2] <= result_col59[1];
   result_col59[3] <= result_col59[2];
   result_col59[4] <= result_col59[3];
   result_col59[5] <= result_col59[4];
   result_col59[6] <= result_col59[5];
   result_col59[7] <= result_col59[6];
   result_col59[8] <= result_col59[7];
   result_col59[9] <= result_col59[8];
   result_col59[10] <= result_col59[9];
   result_col59[11] <= result_col59[10];
   result_col59[12] <= result_col59[11];
   result_col59[13] <= result_col59[12];
   result_col59[14] <= result_col59[13];
   result_col59[15] <= result_col59[14];
   result_col59[16] <= result_col59[15];
   result_col59[17] <= result_col59[16];
   result_col59[18] <= result_col59[17];
   result_col59[19] <= result_col59[18];
   result_col59[20] <= result_col59[19];
   result_col59[21] <= result_col59[20];
   result_col59[22] <= result_col59[21];
   result_col59[23] <= result_col59[22];
   result_col59[24] <= result_col59[23];
   result_col59[25] <= result_col59[24];
   result_col59[26] <= result_col59[25];
   result_col59[27] <= result_col59[26];
   result_col59[28] <= result_col59[27];
   result_col59[29] <= result_col59[28];
   result_col59[30] <= result_col59[29];
   result_col59[31] <= result_col59[30];
   result_col59[32] <= result_col59[31];
   result_col59[33] <= result_col59[32];
   result_col59[34] <= result_col59[33];
   result_col59[35] <= result_col59[34];
   result_col59[36] <= result_col59[35];
   result_col59[37] <= result_col59[36];
   result_col59[38] <= result_col59[37];
   result_col59[39] <= result_col59[38];
   result_col59[40] <= result_col59[39];
   result_col59[41] <= result_col59[40];

   result_col60[1] <= data_out_5_60;
   result_col60[2] <= result_col60[1];
   result_col60[3] <= result_col60[2];
   result_col60[4] <= result_col60[3];
   result_col60[5] <= result_col60[4];
   result_col60[6] <= result_col60[5];
   result_col60[7] <= result_col60[6];
   result_col60[8] <= result_col60[7];
   result_col60[9] <= result_col60[8];
   result_col60[10] <= result_col60[9];
   result_col60[11] <= result_col60[10];
   result_col60[12] <= result_col60[11];
   result_col60[13] <= result_col60[12];
   result_col60[14] <= result_col60[13];
   result_col60[15] <= result_col60[14];
   result_col60[16] <= result_col60[15];
   result_col60[17] <= result_col60[16];
   result_col60[18] <= result_col60[17];
   result_col60[19] <= result_col60[18];
   result_col60[20] <= result_col60[19];
   result_col60[21] <= result_col60[20];
   result_col60[22] <= result_col60[21];
   result_col60[23] <= result_col60[22];
   result_col60[24] <= result_col60[23];
   result_col60[25] <= result_col60[24];
   result_col60[26] <= result_col60[25];
   result_col60[27] <= result_col60[26];
   result_col60[28] <= result_col60[27];
   result_col60[29] <= result_col60[28];
   result_col60[30] <= result_col60[29];
   result_col60[31] <= result_col60[30];
   result_col60[32] <= result_col60[31];
   result_col60[33] <= result_col60[32];
   result_col60[34] <= result_col60[33];
   result_col60[35] <= result_col60[34];
   result_col60[36] <= result_col60[35];
   result_col60[37] <= result_col60[36];
   result_col60[38] <= result_col60[37];
   result_col60[39] <= result_col60[38];
   result_col60[40] <= result_col60[39];

   result_col61[1] <= data_out_5_61;
   result_col61[2] <= result_col61[1];
   result_col61[3] <= result_col61[2];
   result_col61[4] <= result_col61[3];
   result_col61[5] <= result_col61[4];
   result_col61[6] <= result_col61[5];
   result_col61[7] <= result_col61[6];
   result_col61[8] <= result_col61[7];
   result_col61[9] <= result_col61[8];
   result_col61[10] <= result_col61[9];
   result_col61[11] <= result_col61[10];
   result_col61[12] <= result_col61[11];
   result_col61[13] <= result_col61[12];
   result_col61[14] <= result_col61[13];
   result_col61[15] <= result_col61[14];
   result_col61[16] <= result_col61[15];
   result_col61[17] <= result_col61[16];
   result_col61[18] <= result_col61[17];
   result_col61[19] <= result_col61[18];
   result_col61[20] <= result_col61[19];
   result_col61[21] <= result_col61[20];
   result_col61[22] <= result_col61[21];
   result_col61[23] <= result_col61[22];
   result_col61[24] <= result_col61[23];
   result_col61[25] <= result_col61[24];
   result_col61[26] <= result_col61[25];
   result_col61[27] <= result_col61[26];
   result_col61[28] <= result_col61[27];
   result_col61[29] <= result_col61[28];
   result_col61[30] <= result_col61[29];
   result_col61[31] <= result_col61[30];
   result_col61[32] <= result_col61[31];
   result_col61[33] <= result_col61[32];
   result_col61[34] <= result_col61[33];
   result_col61[35] <= result_col61[34];
   result_col61[36] <= result_col61[35];
   result_col61[37] <= result_col61[36];
   result_col61[38] <= result_col61[37];
   result_col61[39] <= result_col61[38];

   result_col62[1] <= data_out_5_62;
   result_col62[2] <= result_col62[1];
   result_col62[3] <= result_col62[2];
   result_col62[4] <= result_col62[3];
   result_col62[5] <= result_col62[4];
   result_col62[6] <= result_col62[5];
   result_col62[7] <= result_col62[6];
   result_col62[8] <= result_col62[7];
   result_col62[9] <= result_col62[8];
   result_col62[10] <= result_col62[9];
   result_col62[11] <= result_col62[10];
   result_col62[12] <= result_col62[11];
   result_col62[13] <= result_col62[12];
   result_col62[14] <= result_col62[13];
   result_col62[15] <= result_col62[14];
   result_col62[16] <= result_col62[15];
   result_col62[17] <= result_col62[16];
   result_col62[18] <= result_col62[17];
   result_col62[19] <= result_col62[18];
   result_col62[20] <= result_col62[19];
   result_col62[21] <= result_col62[20];
   result_col62[22] <= result_col62[21];
   result_col62[23] <= result_col62[22];
   result_col62[24] <= result_col62[23];
   result_col62[25] <= result_col62[24];
   result_col62[26] <= result_col62[25];
   result_col62[27] <= result_col62[26];
   result_col62[28] <= result_col62[27];
   result_col62[29] <= result_col62[28];
   result_col62[30] <= result_col62[29];
   result_col62[31] <= result_col62[30];
   result_col62[32] <= result_col62[31];
   result_col62[33] <= result_col62[32];
   result_col62[34] <= result_col62[33];
   result_col62[35] <= result_col62[34];
   result_col62[36] <= result_col62[35];
   result_col62[37] <= result_col62[36];
   result_col62[38] <= result_col62[37];

   result_col63[1] <= data_out_5_63;
   result_col63[2] <= result_col63[1];
   result_col63[3] <= result_col63[2];
   result_col63[4] <= result_col63[3];
   result_col63[5] <= result_col63[4];
   result_col63[6] <= result_col63[5];
   result_col63[7] <= result_col63[6];
   result_col63[8] <= result_col63[7];
   result_col63[9] <= result_col63[8];
   result_col63[10] <= result_col63[9];
   result_col63[11] <= result_col63[10];
   result_col63[12] <= result_col63[11];
   result_col63[13] <= result_col63[12];
   result_col63[14] <= result_col63[13];
   result_col63[15] <= result_col63[14];
   result_col63[16] <= result_col63[15];
   result_col63[17] <= result_col63[16];
   result_col63[18] <= result_col63[17];
   result_col63[19] <= result_col63[18];
   result_col63[20] <= result_col63[19];
   result_col63[21] <= result_col63[20];
   result_col63[22] <= result_col63[21];
   result_col63[23] <= result_col63[22];
   result_col63[24] <= result_col63[23];
   result_col63[25] <= result_col63[24];
   result_col63[26] <= result_col63[25];
   result_col63[27] <= result_col63[26];
   result_col63[28] <= result_col63[27];
   result_col63[29] <= result_col63[28];
   result_col63[30] <= result_col63[29];
   result_col63[31] <= result_col63[30];
   result_col63[32] <= result_col63[31];
   result_col63[33] <= result_col63[32];
   result_col63[34] <= result_col63[33];
   result_col63[35] <= result_col63[34];
   result_col63[36] <= result_col63[35];
   result_col63[37] <= result_col63[36];

   result_col64[1] <= data_out_5_64;
   result_col64[2] <= result_col64[1];
   result_col64[3] <= result_col64[2];
   result_col64[4] <= result_col64[3];
   result_col64[5] <= result_col64[4];
   result_col64[6] <= result_col64[5];
   result_col64[7] <= result_col64[6];
   result_col64[8] <= result_col64[7];
   result_col64[9] <= result_col64[8];
   result_col64[10] <= result_col64[9];
   result_col64[11] <= result_col64[10];
   result_col64[12] <= result_col64[11];
   result_col64[13] <= result_col64[12];
   result_col64[14] <= result_col64[13];
   result_col64[15] <= result_col64[14];
   result_col64[16] <= result_col64[15];
   result_col64[17] <= result_col64[16];
   result_col64[18] <= result_col64[17];
   result_col64[19] <= result_col64[18];
   result_col64[20] <= result_col64[19];
   result_col64[21] <= result_col64[20];
   result_col64[22] <= result_col64[21];
   result_col64[23] <= result_col64[22];
   result_col64[24] <= result_col64[23];
   result_col64[25] <= result_col64[24];
   result_col64[26] <= result_col64[25];
   result_col64[27] <= result_col64[26];
   result_col64[28] <= result_col64[27];
   result_col64[29] <= result_col64[28];
   result_col64[30] <= result_col64[29];
   result_col64[31] <= result_col64[30];
   result_col64[32] <= result_col64[31];
   result_col64[33] <= result_col64[32];
   result_col64[34] <= result_col64[33];
   result_col64[35] <= result_col64[34];
   result_col64[36] <= result_col64[35];

   result_col65[1] <= data_out_5_65;
   result_col65[2] <= result_col65[1];
   result_col65[3] <= result_col65[2];
   result_col65[4] <= result_col65[3];
   result_col65[5] <= result_col65[4];
   result_col65[6] <= result_col65[5];
   result_col65[7] <= result_col65[6];
   result_col65[8] <= result_col65[7];
   result_col65[9] <= result_col65[8];
   result_col65[10] <= result_col65[9];
   result_col65[11] <= result_col65[10];
   result_col65[12] <= result_col65[11];
   result_col65[13] <= result_col65[12];
   result_col65[14] <= result_col65[13];
   result_col65[15] <= result_col65[14];
   result_col65[16] <= result_col65[15];
   result_col65[17] <= result_col65[16];
   result_col65[18] <= result_col65[17];
   result_col65[19] <= result_col65[18];
   result_col65[20] <= result_col65[19];
   result_col65[21] <= result_col65[20];
   result_col65[22] <= result_col65[21];
   result_col65[23] <= result_col65[22];
   result_col65[24] <= result_col65[23];
   result_col65[25] <= result_col65[24];
   result_col65[26] <= result_col65[25];
   result_col65[27] <= result_col65[26];
   result_col65[28] <= result_col65[27];
   result_col65[29] <= result_col65[28];
   result_col65[30] <= result_col65[29];
   result_col65[31] <= result_col65[30];
   result_col65[32] <= result_col65[31];
   result_col65[33] <= result_col65[32];
   result_col65[34] <= result_col65[33];
   result_col65[35] <= result_col65[34];

   result_col66[1] <= data_out_5_66;
   result_col66[2] <= result_col66[1];
   result_col66[3] <= result_col66[2];
   result_col66[4] <= result_col66[3];
   result_col66[5] <= result_col66[4];
   result_col66[6] <= result_col66[5];
   result_col66[7] <= result_col66[6];
   result_col66[8] <= result_col66[7];
   result_col66[9] <= result_col66[8];
   result_col66[10] <= result_col66[9];
   result_col66[11] <= result_col66[10];
   result_col66[12] <= result_col66[11];
   result_col66[13] <= result_col66[12];
   result_col66[14] <= result_col66[13];
   result_col66[15] <= result_col66[14];
   result_col66[16] <= result_col66[15];
   result_col66[17] <= result_col66[16];
   result_col66[18] <= result_col66[17];
   result_col66[19] <= result_col66[18];
   result_col66[20] <= result_col66[19];
   result_col66[21] <= result_col66[20];
   result_col66[22] <= result_col66[21];
   result_col66[23] <= result_col66[22];
   result_col66[24] <= result_col66[23];
   result_col66[25] <= result_col66[24];
   result_col66[26] <= result_col66[25];
   result_col66[27] <= result_col66[26];
   result_col66[28] <= result_col66[27];
   result_col66[29] <= result_col66[28];
   result_col66[30] <= result_col66[29];
   result_col66[31] <= result_col66[30];
   result_col66[32] <= result_col66[31];
   result_col66[33] <= result_col66[32];
   result_col66[34] <= result_col66[33];

   result_col67[1] <= data_out_5_67;
   result_col67[2] <= result_col67[1];
   result_col67[3] <= result_col67[2];
   result_col67[4] <= result_col67[3];
   result_col67[5] <= result_col67[4];
   result_col67[6] <= result_col67[5];
   result_col67[7] <= result_col67[6];
   result_col67[8] <= result_col67[7];
   result_col67[9] <= result_col67[8];
   result_col67[10] <= result_col67[9];
   result_col67[11] <= result_col67[10];
   result_col67[12] <= result_col67[11];
   result_col67[13] <= result_col67[12];
   result_col67[14] <= result_col67[13];
   result_col67[15] <= result_col67[14];
   result_col67[16] <= result_col67[15];
   result_col67[17] <= result_col67[16];
   result_col67[18] <= result_col67[17];
   result_col67[19] <= result_col67[18];
   result_col67[20] <= result_col67[19];
   result_col67[21] <= result_col67[20];
   result_col67[22] <= result_col67[21];
   result_col67[23] <= result_col67[22];
   result_col67[24] <= result_col67[23];
   result_col67[25] <= result_col67[24];
   result_col67[26] <= result_col67[25];
   result_col67[27] <= result_col67[26];
   result_col67[28] <= result_col67[27];
   result_col67[29] <= result_col67[28];
   result_col67[30] <= result_col67[29];
   result_col67[31] <= result_col67[30];
   result_col67[32] <= result_col67[31];
   result_col67[33] <= result_col67[32];

   result_col68[1] <= data_out_5_68;
   result_col68[2] <= result_col68[1];
   result_col68[3] <= result_col68[2];
   result_col68[4] <= result_col68[3];
   result_col68[5] <= result_col68[4];
   result_col68[6] <= result_col68[5];
   result_col68[7] <= result_col68[6];
   result_col68[8] <= result_col68[7];
   result_col68[9] <= result_col68[8];
   result_col68[10] <= result_col68[9];
   result_col68[11] <= result_col68[10];
   result_col68[12] <= result_col68[11];
   result_col68[13] <= result_col68[12];
   result_col68[14] <= result_col68[13];
   result_col68[15] <= result_col68[14];
   result_col68[16] <= result_col68[15];
   result_col68[17] <= result_col68[16];
   result_col68[18] <= result_col68[17];
   result_col68[19] <= result_col68[18];
   result_col68[20] <= result_col68[19];
   result_col68[21] <= result_col68[20];
   result_col68[22] <= result_col68[21];
   result_col68[23] <= result_col68[22];
   result_col68[24] <= result_col68[23];
   result_col68[25] <= result_col68[24];
   result_col68[26] <= result_col68[25];
   result_col68[27] <= result_col68[26];
   result_col68[28] <= result_col68[27];
   result_col68[29] <= result_col68[28];
   result_col68[30] <= result_col68[29];
   result_col68[31] <= result_col68[30];
   result_col68[32] <= result_col68[31];

   result_col69[1] <= data_out_5_69;
   result_col69[2] <= result_col69[1];
   result_col69[3] <= result_col69[2];
   result_col69[4] <= result_col69[3];
   result_col69[5] <= result_col69[4];
   result_col69[6] <= result_col69[5];
   result_col69[7] <= result_col69[6];
   result_col69[8] <= result_col69[7];
   result_col69[9] <= result_col69[8];
   result_col69[10] <= result_col69[9];
   result_col69[11] <= result_col69[10];
   result_col69[12] <= result_col69[11];
   result_col69[13] <= result_col69[12];
   result_col69[14] <= result_col69[13];
   result_col69[15] <= result_col69[14];
   result_col69[16] <= result_col69[15];
   result_col69[17] <= result_col69[16];
   result_col69[18] <= result_col69[17];
   result_col69[19] <= result_col69[18];
   result_col69[20] <= result_col69[19];
   result_col69[21] <= result_col69[20];
   result_col69[22] <= result_col69[21];
   result_col69[23] <= result_col69[22];
   result_col69[24] <= result_col69[23];
   result_col69[25] <= result_col69[24];
   result_col69[26] <= result_col69[25];
   result_col69[27] <= result_col69[26];
   result_col69[28] <= result_col69[27];
   result_col69[29] <= result_col69[28];
   result_col69[30] <= result_col69[29];
   result_col69[31] <= result_col69[30];

   result_col70[1] <= data_out_5_70;
   result_col70[2] <= result_col70[1];
   result_col70[3] <= result_col70[2];
   result_col70[4] <= result_col70[3];
   result_col70[5] <= result_col70[4];
   result_col70[6] <= result_col70[5];
   result_col70[7] <= result_col70[6];
   result_col70[8] <= result_col70[7];
   result_col70[9] <= result_col70[8];
   result_col70[10] <= result_col70[9];
   result_col70[11] <= result_col70[10];
   result_col70[12] <= result_col70[11];
   result_col70[13] <= result_col70[12];
   result_col70[14] <= result_col70[13];
   result_col70[15] <= result_col70[14];
   result_col70[16] <= result_col70[15];
   result_col70[17] <= result_col70[16];
   result_col70[18] <= result_col70[17];
   result_col70[19] <= result_col70[18];
   result_col70[20] <= result_col70[19];
   result_col70[21] <= result_col70[20];
   result_col70[22] <= result_col70[21];
   result_col70[23] <= result_col70[22];
   result_col70[24] <= result_col70[23];
   result_col70[25] <= result_col70[24];
   result_col70[26] <= result_col70[25];
   result_col70[27] <= result_col70[26];
   result_col70[28] <= result_col70[27];
   result_col70[29] <= result_col70[28];
   result_col70[30] <= result_col70[29];

   result_col71[1] <= data_out_5_71;
   result_col71[2] <= result_col71[1];
   result_col71[3] <= result_col71[2];
   result_col71[4] <= result_col71[3];
   result_col71[5] <= result_col71[4];
   result_col71[6] <= result_col71[5];
   result_col71[7] <= result_col71[6];
   result_col71[8] <= result_col71[7];
   result_col71[9] <= result_col71[8];
   result_col71[10] <= result_col71[9];
   result_col71[11] <= result_col71[10];
   result_col71[12] <= result_col71[11];
   result_col71[13] <= result_col71[12];
   result_col71[14] <= result_col71[13];
   result_col71[15] <= result_col71[14];
   result_col71[16] <= result_col71[15];
   result_col71[17] <= result_col71[16];
   result_col71[18] <= result_col71[17];
   result_col71[19] <= result_col71[18];
   result_col71[20] <= result_col71[19];
   result_col71[21] <= result_col71[20];
   result_col71[22] <= result_col71[21];
   result_col71[23] <= result_col71[22];
   result_col71[24] <= result_col71[23];
   result_col71[25] <= result_col71[24];
   result_col71[26] <= result_col71[25];
   result_col71[27] <= result_col71[26];
   result_col71[28] <= result_col71[27];
   result_col71[29] <= result_col71[28];

   result_col72[1] <= data_out_5_72;
   result_col72[2] <= result_col72[1];
   result_col72[3] <= result_col72[2];
   result_col72[4] <= result_col72[3];
   result_col72[5] <= result_col72[4];
   result_col72[6] <= result_col72[5];
   result_col72[7] <= result_col72[6];
   result_col72[8] <= result_col72[7];
   result_col72[9] <= result_col72[8];
   result_col72[10] <= result_col72[9];
   result_col72[11] <= result_col72[10];
   result_col72[12] <= result_col72[11];
   result_col72[13] <= result_col72[12];
   result_col72[14] <= result_col72[13];
   result_col72[15] <= result_col72[14];
   result_col72[16] <= result_col72[15];
   result_col72[17] <= result_col72[16];
   result_col72[18] <= result_col72[17];
   result_col72[19] <= result_col72[18];
   result_col72[20] <= result_col72[19];
   result_col72[21] <= result_col72[20];
   result_col72[22] <= result_col72[21];
   result_col72[23] <= result_col72[22];
   result_col72[24] <= result_col72[23];
   result_col72[25] <= result_col72[24];
   result_col72[26] <= result_col72[25];
   result_col72[27] <= result_col72[26];
   result_col72[28] <= result_col72[27];

   result_col73[1] <= data_out_5_73;
   result_col73[2] <= result_col73[1];
   result_col73[3] <= result_col73[2];
   result_col73[4] <= result_col73[3];
   result_col73[5] <= result_col73[4];
   result_col73[6] <= result_col73[5];
   result_col73[7] <= result_col73[6];
   result_col73[8] <= result_col73[7];
   result_col73[9] <= result_col73[8];
   result_col73[10] <= result_col73[9];
   result_col73[11] <= result_col73[10];
   result_col73[12] <= result_col73[11];
   result_col73[13] <= result_col73[12];
   result_col73[14] <= result_col73[13];
   result_col73[15] <= result_col73[14];
   result_col73[16] <= result_col73[15];
   result_col73[17] <= result_col73[16];
   result_col73[18] <= result_col73[17];
   result_col73[19] <= result_col73[18];
   result_col73[20] <= result_col73[19];
   result_col73[21] <= result_col73[20];
   result_col73[22] <= result_col73[21];
   result_col73[23] <= result_col73[22];
   result_col73[24] <= result_col73[23];
   result_col73[25] <= result_col73[24];
   result_col73[26] <= result_col73[25];
   result_col73[27] <= result_col73[26];

   result_col74[1] <= data_out_5_74;
   result_col74[2] <= result_col74[1];
   result_col74[3] <= result_col74[2];
   result_col74[4] <= result_col74[3];
   result_col74[5] <= result_col74[4];
   result_col74[6] <= result_col74[5];
   result_col74[7] <= result_col74[6];
   result_col74[8] <= result_col74[7];
   result_col74[9] <= result_col74[8];
   result_col74[10] <= result_col74[9];
   result_col74[11] <= result_col74[10];
   result_col74[12] <= result_col74[11];
   result_col74[13] <= result_col74[12];
   result_col74[14] <= result_col74[13];
   result_col74[15] <= result_col74[14];
   result_col74[16] <= result_col74[15];
   result_col74[17] <= result_col74[16];
   result_col74[18] <= result_col74[17];
   result_col74[19] <= result_col74[18];
   result_col74[20] <= result_col74[19];
   result_col74[21] <= result_col74[20];
   result_col74[22] <= result_col74[21];
   result_col74[23] <= result_col74[22];
   result_col74[24] <= result_col74[23];
   result_col74[25] <= result_col74[24];
   result_col74[26] <= result_col74[25];

   result_col75[1] <= data_out_5_75;
   result_col75[2] <= result_col75[1];
   result_col75[3] <= result_col75[2];
   result_col75[4] <= result_col75[3];
   result_col75[5] <= result_col75[4];
   result_col75[6] <= result_col75[5];
   result_col75[7] <= result_col75[6];
   result_col75[8] <= result_col75[7];
   result_col75[9] <= result_col75[8];
   result_col75[10] <= result_col75[9];
   result_col75[11] <= result_col75[10];
   result_col75[12] <= result_col75[11];
   result_col75[13] <= result_col75[12];
   result_col75[14] <= result_col75[13];
   result_col75[15] <= result_col75[14];
   result_col75[16] <= result_col75[15];
   result_col75[17] <= result_col75[16];
   result_col75[18] <= result_col75[17];
   result_col75[19] <= result_col75[18];
   result_col75[20] <= result_col75[19];
   result_col75[21] <= result_col75[20];
   result_col75[22] <= result_col75[21];
   result_col75[23] <= result_col75[22];
   result_col75[24] <= result_col75[23];
   result_col75[25] <= result_col75[24];

   result_col76[1] <= data_out_5_76;
   result_col76[2] <= result_col76[1];
   result_col76[3] <= result_col76[2];
   result_col76[4] <= result_col76[3];
   result_col76[5] <= result_col76[4];
   result_col76[6] <= result_col76[5];
   result_col76[7] <= result_col76[6];
   result_col76[8] <= result_col76[7];
   result_col76[9] <= result_col76[8];
   result_col76[10] <= result_col76[9];
   result_col76[11] <= result_col76[10];
   result_col76[12] <= result_col76[11];
   result_col76[13] <= result_col76[12];
   result_col76[14] <= result_col76[13];
   result_col76[15] <= result_col76[14];
   result_col76[16] <= result_col76[15];
   result_col76[17] <= result_col76[16];
   result_col76[18] <= result_col76[17];
   result_col76[19] <= result_col76[18];
   result_col76[20] <= result_col76[19];
   result_col76[21] <= result_col76[20];
   result_col76[22] <= result_col76[21];
   result_col76[23] <= result_col76[22];
   result_col76[24] <= result_col76[23];

   result_col77[1] <= data_out_5_77;
   result_col77[2] <= result_col77[1];
   result_col77[3] <= result_col77[2];
   result_col77[4] <= result_col77[3];
   result_col77[5] <= result_col77[4];
   result_col77[6] <= result_col77[5];
   result_col77[7] <= result_col77[6];
   result_col77[8] <= result_col77[7];
   result_col77[9] <= result_col77[8];
   result_col77[10] <= result_col77[9];
   result_col77[11] <= result_col77[10];
   result_col77[12] <= result_col77[11];
   result_col77[13] <= result_col77[12];
   result_col77[14] <= result_col77[13];
   result_col77[15] <= result_col77[14];
   result_col77[16] <= result_col77[15];
   result_col77[17] <= result_col77[16];
   result_col77[18] <= result_col77[17];
   result_col77[19] <= result_col77[18];
   result_col77[20] <= result_col77[19];
   result_col77[21] <= result_col77[20];
   result_col77[22] <= result_col77[21];
   result_col77[23] <= result_col77[22];

   result_col78[1] <= data_out_5_78;
   result_col78[2] <= result_col78[1];
   result_col78[3] <= result_col78[2];
   result_col78[4] <= result_col78[3];
   result_col78[5] <= result_col78[4];
   result_col78[6] <= result_col78[5];
   result_col78[7] <= result_col78[6];
   result_col78[8] <= result_col78[7];
   result_col78[9] <= result_col78[8];
   result_col78[10] <= result_col78[9];
   result_col78[11] <= result_col78[10];
   result_col78[12] <= result_col78[11];
   result_col78[13] <= result_col78[12];
   result_col78[14] <= result_col78[13];
   result_col78[15] <= result_col78[14];
   result_col78[16] <= result_col78[15];
   result_col78[17] <= result_col78[16];
   result_col78[18] <= result_col78[17];
   result_col78[19] <= result_col78[18];
   result_col78[20] <= result_col78[19];
   result_col78[21] <= result_col78[20];
   result_col78[22] <= result_col78[21];

   result_col79[1] <= data_out_5_79;
   result_col79[2] <= result_col79[1];
   result_col79[3] <= result_col79[2];
   result_col79[4] <= result_col79[3];
   result_col79[5] <= result_col79[4];
   result_col79[6] <= result_col79[5];
   result_col79[7] <= result_col79[6];
   result_col79[8] <= result_col79[7];
   result_col79[9] <= result_col79[8];
   result_col79[10] <= result_col79[9];
   result_col79[11] <= result_col79[10];
   result_col79[12] <= result_col79[11];
   result_col79[13] <= result_col79[12];
   result_col79[14] <= result_col79[13];
   result_col79[15] <= result_col79[14];
   result_col79[16] <= result_col79[15];
   result_col79[17] <= result_col79[16];
   result_col79[18] <= result_col79[17];
   result_col79[19] <= result_col79[18];
   result_col79[20] <= result_col79[19];
   result_col79[21] <= result_col79[20];

   result_col80[1] <= data_out_5_80;
   result_col80[2] <= result_col80[1];
   result_col80[3] <= result_col80[2];
   result_col80[4] <= result_col80[3];
   result_col80[5] <= result_col80[4];
   result_col80[6] <= result_col80[5];
   result_col80[7] <= result_col80[6];
   result_col80[8] <= result_col80[7];
   result_col80[9] <= result_col80[8];
   result_col80[10] <= result_col80[9];
   result_col80[11] <= result_col80[10];
   result_col80[12] <= result_col80[11];
   result_col80[13] <= result_col80[12];
   result_col80[14] <= result_col80[13];
   result_col80[15] <= result_col80[14];
   result_col80[16] <= result_col80[15];
   result_col80[17] <= result_col80[16];
   result_col80[18] <= result_col80[17];
   result_col80[19] <= result_col80[18];
   result_col80[20] <= result_col80[19];

   result_col81[1] <= data_out_5_81;
   result_col81[2] <= result_col81[1];
   result_col81[3] <= result_col81[2];
   result_col81[4] <= result_col81[3];
   result_col81[5] <= result_col81[4];
   result_col81[6] <= result_col81[5];
   result_col81[7] <= result_col81[6];
   result_col81[8] <= result_col81[7];
   result_col81[9] <= result_col81[8];
   result_col81[10] <= result_col81[9];
   result_col81[11] <= result_col81[10];
   result_col81[12] <= result_col81[11];
   result_col81[13] <= result_col81[12];
   result_col81[14] <= result_col81[13];
   result_col81[15] <= result_col81[14];
   result_col81[16] <= result_col81[15];
   result_col81[17] <= result_col81[16];
   result_col81[18] <= result_col81[17];
   result_col81[19] <= result_col81[18];

   result_col82[1] <= data_out_5_82;
   result_col82[2] <= result_col82[1];
   result_col82[3] <= result_col82[2];
   result_col82[4] <= result_col82[3];
   result_col82[5] <= result_col82[4];
   result_col82[6] <= result_col82[5];
   result_col82[7] <= result_col82[6];
   result_col82[8] <= result_col82[7];
   result_col82[9] <= result_col82[8];
   result_col82[10] <= result_col82[9];
   result_col82[11] <= result_col82[10];
   result_col82[12] <= result_col82[11];
   result_col82[13] <= result_col82[12];
   result_col82[14] <= result_col82[13];
   result_col82[15] <= result_col82[14];
   result_col82[16] <= result_col82[15];
   result_col82[17] <= result_col82[16];
   result_col82[18] <= result_col82[17];

   result_col83[1] <= data_out_5_83;
   result_col83[2] <= result_col83[1];
   result_col83[3] <= result_col83[2];
   result_col83[4] <= result_col83[3];
   result_col83[5] <= result_col83[4];
   result_col83[6] <= result_col83[5];
   result_col83[7] <= result_col83[6];
   result_col83[8] <= result_col83[7];
   result_col83[9] <= result_col83[8];
   result_col83[10] <= result_col83[9];
   result_col83[11] <= result_col83[10];
   result_col83[12] <= result_col83[11];
   result_col83[13] <= result_col83[12];
   result_col83[14] <= result_col83[13];
   result_col83[15] <= result_col83[14];
   result_col83[16] <= result_col83[15];
   result_col83[17] <= result_col83[16];

   result_col84[1] <= data_out_5_84;
   result_col84[2] <= result_col84[1];
   result_col84[3] <= result_col84[2];
   result_col84[4] <= result_col84[3];
   result_col84[5] <= result_col84[4];
   result_col84[6] <= result_col84[5];
   result_col84[7] <= result_col84[6];
   result_col84[8] <= result_col84[7];
   result_col84[9] <= result_col84[8];
   result_col84[10] <= result_col84[9];
   result_col84[11] <= result_col84[10];
   result_col84[12] <= result_col84[11];
   result_col84[13] <= result_col84[12];
   result_col84[14] <= result_col84[13];
   result_col84[15] <= result_col84[14];
   result_col84[16] <= result_col84[15];

   result_col85[1] <= data_out_5_85;
   result_col85[2] <= result_col85[1];
   result_col85[3] <= result_col85[2];
   result_col85[4] <= result_col85[3];
   result_col85[5] <= result_col85[4];
   result_col85[6] <= result_col85[5];
   result_col85[7] <= result_col85[6];
   result_col85[8] <= result_col85[7];
   result_col85[9] <= result_col85[8];
   result_col85[10] <= result_col85[9];
   result_col85[11] <= result_col85[10];
   result_col85[12] <= result_col85[11];
   result_col85[13] <= result_col85[12];
   result_col85[14] <= result_col85[13];
   result_col85[15] <= result_col85[14];

   result_col86[1] <= data_out_5_86;
   result_col86[2] <= result_col86[1];
   result_col86[3] <= result_col86[2];
   result_col86[4] <= result_col86[3];
   result_col86[5] <= result_col86[4];
   result_col86[6] <= result_col86[5];
   result_col86[7] <= result_col86[6];
   result_col86[8] <= result_col86[7];
   result_col86[9] <= result_col86[8];
   result_col86[10] <= result_col86[9];
   result_col86[11] <= result_col86[10];
   result_col86[12] <= result_col86[11];
   result_col86[13] <= result_col86[12];
   result_col86[14] <= result_col86[13];

   result_col87[1] <= data_out_5_87;
   result_col87[2] <= result_col87[1];
   result_col87[3] <= result_col87[2];
   result_col87[4] <= result_col87[3];
   result_col87[5] <= result_col87[4];
   result_col87[6] <= result_col87[5];
   result_col87[7] <= result_col87[6];
   result_col87[8] <= result_col87[7];
   result_col87[9] <= result_col87[8];
   result_col87[10] <= result_col87[9];
   result_col87[11] <= result_col87[10];
   result_col87[12] <= result_col87[11];
   result_col87[13] <= result_col87[12];

   result_col88[1] <= data_out_5_88;
   result_col88[2] <= result_col88[1];
   result_col88[3] <= result_col88[2];
   result_col88[4] <= result_col88[3];
   result_col88[5] <= result_col88[4];
   result_col88[6] <= result_col88[5];
   result_col88[7] <= result_col88[6];
   result_col88[8] <= result_col88[7];
   result_col88[9] <= result_col88[8];
   result_col88[10] <= result_col88[9];
   result_col88[11] <= result_col88[10];
   result_col88[12] <= result_col88[11];

   result_col89[1] <= data_out_5_89;
   result_col89[2] <= result_col89[1];
   result_col89[3] <= result_col89[2];
   result_col89[4] <= result_col89[3];
   result_col89[5] <= result_col89[4];
   result_col89[6] <= result_col89[5];
   result_col89[7] <= result_col89[6];
   result_col89[8] <= result_col89[7];
   result_col89[9] <= result_col89[8];
   result_col89[10] <= result_col89[9];
   result_col89[11] <= result_col89[10];

   result_col90[1] <= data_out_5_90;
   result_col90[2] <= result_col90[1];
   result_col90[3] <= result_col90[2];
   result_col90[4] <= result_col90[3];
   result_col90[5] <= result_col90[4];
   result_col90[6] <= result_col90[5];
   result_col90[7] <= result_col90[6];
   result_col90[8] <= result_col90[7];
   result_col90[9] <= result_col90[8];
   result_col90[10] <= result_col90[9];

   result_col91[1] <= data_out_5_91;
   result_col91[2] <= result_col91[1];
   result_col91[3] <= result_col91[2];
   result_col91[4] <= result_col91[3];
   result_col91[5] <= result_col91[4];
   result_col91[6] <= result_col91[5];
   result_col91[7] <= result_col91[6];
   result_col91[8] <= result_col91[7];
   result_col91[9] <= result_col91[8];

   result_col92[1] <= data_out_5_92;
   result_col92[2] <= result_col92[1];
   result_col92[3] <= result_col92[2];
   result_col92[4] <= result_col92[3];
   result_col92[5] <= result_col92[4];
   result_col92[6] <= result_col92[5];
   result_col92[7] <= result_col92[6];
   result_col92[8] <= result_col92[7];

   result_col93[1] <= data_out_5_93;
   result_col93[2] <= result_col93[1];
   result_col93[3] <= result_col93[2];
   result_col93[4] <= result_col93[3];
   result_col93[5] <= result_col93[4];
   result_col93[6] <= result_col93[5];
   result_col93[7] <= result_col93[6];

   result_col94[1] <= data_out_5_94;
   result_col94[2] <= result_col94[1];
   result_col94[3] <= result_col94[2];
   result_col94[4] <= result_col94[3];
   result_col94[5] <= result_col94[4];
   result_col94[6] <= result_col94[5];

   result_col95[1] <= data_out_5_95;
   result_col95[2] <= result_col95[1];
   result_col95[3] <= result_col95[2];
   result_col95[4] <= result_col95[3];
   result_col95[5] <= result_col95[4];

   result_col96[1] <= data_out_5_96;
   result_col96[2] <= result_col96[1];
   result_col96[3] <= result_col96[2];
   result_col96[4] <= result_col96[3];

   result_col97[1] <= data_out_5_97;
   result_col97[2] <= result_col97[1];
   result_col97[3] <= result_col97[2];

   result_col98[1] <= data_out_5_98;
   result_col98[2] <= result_col98[1];

   result_col99[1] <= data_out_5_99;
 end

 assign result = {result_col0[100], result_col1[99], result_col2[98], result_col3[97], result_col4[96], result_col5[95], result_col6[94], result_col7[93], result_col8[92], result_col9[91], result_col10[90], result_col11[89], result_col12[88], result_col13[87], result_col14[86], result_col15[85], result_col16[84], result_col17[83], result_col18[82], result_col19[81], result_col20[80], result_col21[79], result_col22[78], result_col23[77], result_col24[76], result_col25[75], result_col26[74], result_col27[73], result_col28[72], result_col29[71], result_col30[70], result_col31[69], result_col32[68], result_col33[67], result_col34[66], result_col35[65], result_col36[64], result_col37[63], result_col38[62], result_col39[61], result_col40[60], result_col41[59], result_col42[58], result_col43[57], result_col44[56], result_col45[55], result_col46[54], result_col47[53], result_col48[52], result_col49[51], result_col50[50], result_col51[49], result_col52[48], result_col53[47], result_col54[46], result_col55[45], result_col56[44], result_col57[43], result_col58[42], result_col59[41], result_col60[40], result_col61[39], result_col62[38], result_col63[37], result_col64[36], result_col65[35], result_col66[34], result_col67[33], result_col68[32], result_col69[31], result_col70[30], result_col71[29], result_col72[28], result_col73[27], result_col74[26], result_col75[25], result_col76[24], result_col77[23], result_col78[22], result_col79[21], result_col80[20], result_col81[19], result_col82[18], result_col83[17], result_col84[16], result_col85[15], result_col86[14], result_col87[13], result_col88[12], result_col89[11], result_col90[10], result_col91[9], result_col92[8], result_col93[7], result_col94[6], result_col95[5], result_col96[4], result_col97[3], result_col98[2], result_col99[1], result_col100};

endmodule

