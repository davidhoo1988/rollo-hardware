module comb_SA #(parameter DAT_W = 166)(
  input wire clk,
  input wire rst_b,
  input wire mode,
  input start,
  input swap,
  input wire [DAT_W-1:0] data,
  output reg finish,
  output wire full_rank,
  output wire [DAT_W-1:0] result
);

  reg [4 : 1] start_tmp;
  reg [4 : 1] start_row;

  reg [4 : 1] swap_row;

  always @(posedge clk) begin
    start_tmp[1] <= start;
    start_row[1] <= start_tmp[1];
    start_tmp[2] <= start_row[1];
    start_row[2] <= start_tmp[2];
    start_tmp[3] <= start_row[2];
    start_row[3] <= start_tmp[3];
    start_tmp[4] <= start_row[3];
    start_row[4] <= start_tmp[4];
  end

  always @(posedge clk) begin
    swap_row[1] <= swap;
    swap_row[2] <= swap_row[1];
    swap_row[3] <= swap_row[2];
    swap_row[4] <= swap_row[3];
  end

 //input skewed form
 wire data_col0;
 reg [1:1] data_col1;
 reg [2:1] data_col2;
 reg [3:1] data_col3;
 reg [4:1] data_col4;
 reg [5:1] data_col5;
 reg [6:1] data_col6;
 reg [7:1] data_col7;
 reg [8:1] data_col8;
 reg [9:1] data_col9;
 reg [10:1] data_col10;
 reg [11:1] data_col11;
 reg [12:1] data_col12;
 reg [13:1] data_col13;
 reg [14:1] data_col14;
 reg [15:1] data_col15;
 reg [16:1] data_col16;
 reg [17:1] data_col17;
 reg [18:1] data_col18;
 reg [19:1] data_col19;
 reg [20:1] data_col20;
 reg [21:1] data_col21;
 reg [22:1] data_col22;
 reg [23:1] data_col23;
 reg [24:1] data_col24;
 reg [25:1] data_col25;
 reg [26:1] data_col26;
 reg [27:1] data_col27;
 reg [28:1] data_col28;
 reg [29:1] data_col29;
 reg [30:1] data_col30;
 reg [31:1] data_col31;
 reg [32:1] data_col32;
 reg [33:1] data_col33;
 reg [34:1] data_col34;
 reg [35:1] data_col35;
 reg [36:1] data_col36;
 reg [37:1] data_col37;
 reg [38:1] data_col38;
 reg [39:1] data_col39;
 reg [40:1] data_col40;
 reg [41:1] data_col41;
 reg [42:1] data_col42;
 reg [43:1] data_col43;
 reg [44:1] data_col44;
 reg [45:1] data_col45;
 reg [46:1] data_col46;
 reg [47:1] data_col47;
 reg [48:1] data_col48;
 reg [49:1] data_col49;
 reg [50:1] data_col50;
 reg [51:1] data_col51;
 reg [52:1] data_col52;
 reg [53:1] data_col53;
 reg [54:1] data_col54;
 reg [55:1] data_col55;
 reg [56:1] data_col56;
 reg [57:1] data_col57;
 reg [58:1] data_col58;
 reg [59:1] data_col59;
 reg [60:1] data_col60;
 reg [61:1] data_col61;
 reg [62:1] data_col62;
 reg [63:1] data_col63;
 reg [64:1] data_col64;
 reg [65:1] data_col65;
 reg [66:1] data_col66;
 reg [67:1] data_col67;
 reg [68:1] data_col68;
 reg [69:1] data_col69;
 reg [70:1] data_col70;
 reg [71:1] data_col71;
 reg [72:1] data_col72;
 reg [73:1] data_col73;
 reg [74:1] data_col74;
 reg [75:1] data_col75;
 reg [76:1] data_col76;
 reg [77:1] data_col77;
 reg [78:1] data_col78;
 reg [79:1] data_col79;
 reg [80:1] data_col80;
 reg [81:1] data_col81;
 reg [82:1] data_col82;
 reg [83:1] data_col83;
 reg [84:1] data_col84;
 reg [85:1] data_col85;
 reg [86:1] data_col86;
 reg [87:1] data_col87;
 reg [88:1] data_col88;
 reg [89:1] data_col89;
 reg [90:1] data_col90;
 reg [91:1] data_col91;
 reg [92:1] data_col92;
 reg [93:1] data_col93;
 reg [94:1] data_col94;
 reg [95:1] data_col95;
 reg [96:1] data_col96;
 reg [97:1] data_col97;
 reg [98:1] data_col98;
 reg [99:1] data_col99;
 reg [100:1] data_col100;
 reg [101:1] data_col101;
 reg [102:1] data_col102;
 reg [103:1] data_col103;
 reg [104:1] data_col104;
 reg [105:1] data_col105;
 reg [106:1] data_col106;
 reg [107:1] data_col107;
 reg [108:1] data_col108;
 reg [109:1] data_col109;
 reg [110:1] data_col110;
 reg [111:1] data_col111;
 reg [112:1] data_col112;
 reg [113:1] data_col113;
 reg [114:1] data_col114;
 reg [115:1] data_col115;
 reg [116:1] data_col116;
 reg [117:1] data_col117;
 reg [118:1] data_col118;
 reg [119:1] data_col119;
 reg [120:1] data_col120;
 reg [121:1] data_col121;
 reg [122:1] data_col122;
 reg [123:1] data_col123;
 reg [124:1] data_col124;
 reg [125:1] data_col125;
 reg [126:1] data_col126;
 reg [127:1] data_col127;
 reg [128:1] data_col128;
 reg [129:1] data_col129;
 reg [130:1] data_col130;
 reg [131:1] data_col131;
 reg [132:1] data_col132;
 reg [133:1] data_col133;
 reg [134:1] data_col134;
 reg [135:1] data_col135;
 reg [136:1] data_col136;
 reg [137:1] data_col137;
 reg [138:1] data_col138;
 reg [139:1] data_col139;
 reg [140:1] data_col140;
 reg [141:1] data_col141;
 reg [142:1] data_col142;
 reg [143:1] data_col143;
 reg [144:1] data_col144;
 reg [145:1] data_col145;
 reg [146:1] data_col146;
 reg [147:1] data_col147;
 reg [148:1] data_col148;
 reg [149:1] data_col149;
 reg [150:1] data_col150;
 reg [151:1] data_col151;
 reg [152:1] data_col152;
 reg [153:1] data_col153;
 reg [154:1] data_col154;
 reg [155:1] data_col155;
 reg [156:1] data_col156;
 reg [157:1] data_col157;
 reg [158:1] data_col158;
 reg [159:1] data_col159;
 reg [160:1] data_col160;
 reg [161:1] data_col161;
 reg [162:1] data_col162;
 reg [163:1] data_col163;
 reg [164:1] data_col164;
 reg [165:1] data_col165;

 assign data_col0 = data[165];

  always @(posedge clk) begin
   data_col1[1] <= data[164];

   data_col2[1] <= data[163];
   data_col2[2] <= data_col2[1];

   data_col3[1] <= data[162];
   data_col3[2] <= data_col3[1];
   data_col3[3] <= data_col3[2];

   data_col4[1] <= data[161];
   data_col4[2] <= data_col4[1];
   data_col4[3] <= data_col4[2];
   data_col4[4] <= data_col4[3];

   data_col5[1] <= data[160];
   data_col5[2] <= data_col5[1];
   data_col5[3] <= data_col5[2];
   data_col5[4] <= data_col5[3];
   data_col5[5] <= data_col5[4];

   data_col6[1] <= data[159];
   data_col6[2] <= data_col6[1];
   data_col6[3] <= data_col6[2];
   data_col6[4] <= data_col6[3];
   data_col6[5] <= data_col6[4];
   data_col6[6] <= data_col6[5];

   data_col7[1] <= data[158];
   data_col7[2] <= data_col7[1];
   data_col7[3] <= data_col7[2];
   data_col7[4] <= data_col7[3];
   data_col7[5] <= data_col7[4];
   data_col7[6] <= data_col7[5];
   data_col7[7] <= data_col7[6];

   data_col8[1] <= data[157];
   data_col8[2] <= data_col8[1];
   data_col8[3] <= data_col8[2];
   data_col8[4] <= data_col8[3];
   data_col8[5] <= data_col8[4];
   data_col8[6] <= data_col8[5];
   data_col8[7] <= data_col8[6];
   data_col8[8] <= data_col8[7];

   data_col9[1] <= data[156];
   data_col9[2] <= data_col9[1];
   data_col9[3] <= data_col9[2];
   data_col9[4] <= data_col9[3];
   data_col9[5] <= data_col9[4];
   data_col9[6] <= data_col9[5];
   data_col9[7] <= data_col9[6];
   data_col9[8] <= data_col9[7];
   data_col9[9] <= data_col9[8];

   data_col10[1] <= data[155];
   data_col10[2] <= data_col10[1];
   data_col10[3] <= data_col10[2];
   data_col10[4] <= data_col10[3];
   data_col10[5] <= data_col10[4];
   data_col10[6] <= data_col10[5];
   data_col10[7] <= data_col10[6];
   data_col10[8] <= data_col10[7];
   data_col10[9] <= data_col10[8];
   data_col10[10] <= data_col10[9];

   data_col11[1] <= data[154];
   data_col11[2] <= data_col11[1];
   data_col11[3] <= data_col11[2];
   data_col11[4] <= data_col11[3];
   data_col11[5] <= data_col11[4];
   data_col11[6] <= data_col11[5];
   data_col11[7] <= data_col11[6];
   data_col11[8] <= data_col11[7];
   data_col11[9] <= data_col11[8];
   data_col11[10] <= data_col11[9];
   data_col11[11] <= data_col11[10];

   data_col12[1] <= data[153];
   data_col12[2] <= data_col12[1];
   data_col12[3] <= data_col12[2];
   data_col12[4] <= data_col12[3];
   data_col12[5] <= data_col12[4];
   data_col12[6] <= data_col12[5];
   data_col12[7] <= data_col12[6];
   data_col12[8] <= data_col12[7];
   data_col12[9] <= data_col12[8];
   data_col12[10] <= data_col12[9];
   data_col12[11] <= data_col12[10];
   data_col12[12] <= data_col12[11];

   data_col13[1] <= data[152];
   data_col13[2] <= data_col13[1];
   data_col13[3] <= data_col13[2];
   data_col13[4] <= data_col13[3];
   data_col13[5] <= data_col13[4];
   data_col13[6] <= data_col13[5];
   data_col13[7] <= data_col13[6];
   data_col13[8] <= data_col13[7];
   data_col13[9] <= data_col13[8];
   data_col13[10] <= data_col13[9];
   data_col13[11] <= data_col13[10];
   data_col13[12] <= data_col13[11];
   data_col13[13] <= data_col13[12];

   data_col14[1] <= data[151];
   data_col14[2] <= data_col14[1];
   data_col14[3] <= data_col14[2];
   data_col14[4] <= data_col14[3];
   data_col14[5] <= data_col14[4];
   data_col14[6] <= data_col14[5];
   data_col14[7] <= data_col14[6];
   data_col14[8] <= data_col14[7];
   data_col14[9] <= data_col14[8];
   data_col14[10] <= data_col14[9];
   data_col14[11] <= data_col14[10];
   data_col14[12] <= data_col14[11];
   data_col14[13] <= data_col14[12];
   data_col14[14] <= data_col14[13];

   data_col15[1] <= data[150];
   data_col15[2] <= data_col15[1];
   data_col15[3] <= data_col15[2];
   data_col15[4] <= data_col15[3];
   data_col15[5] <= data_col15[4];
   data_col15[6] <= data_col15[5];
   data_col15[7] <= data_col15[6];
   data_col15[8] <= data_col15[7];
   data_col15[9] <= data_col15[8];
   data_col15[10] <= data_col15[9];
   data_col15[11] <= data_col15[10];
   data_col15[12] <= data_col15[11];
   data_col15[13] <= data_col15[12];
   data_col15[14] <= data_col15[13];
   data_col15[15] <= data_col15[14];

   data_col16[1] <= data[149];
   data_col16[2] <= data_col16[1];
   data_col16[3] <= data_col16[2];
   data_col16[4] <= data_col16[3];
   data_col16[5] <= data_col16[4];
   data_col16[6] <= data_col16[5];
   data_col16[7] <= data_col16[6];
   data_col16[8] <= data_col16[7];
   data_col16[9] <= data_col16[8];
   data_col16[10] <= data_col16[9];
   data_col16[11] <= data_col16[10];
   data_col16[12] <= data_col16[11];
   data_col16[13] <= data_col16[12];
   data_col16[14] <= data_col16[13];
   data_col16[15] <= data_col16[14];
   data_col16[16] <= data_col16[15];

   data_col17[1] <= data[148];
   data_col17[2] <= data_col17[1];
   data_col17[3] <= data_col17[2];
   data_col17[4] <= data_col17[3];
   data_col17[5] <= data_col17[4];
   data_col17[6] <= data_col17[5];
   data_col17[7] <= data_col17[6];
   data_col17[8] <= data_col17[7];
   data_col17[9] <= data_col17[8];
   data_col17[10] <= data_col17[9];
   data_col17[11] <= data_col17[10];
   data_col17[12] <= data_col17[11];
   data_col17[13] <= data_col17[12];
   data_col17[14] <= data_col17[13];
   data_col17[15] <= data_col17[14];
   data_col17[16] <= data_col17[15];
   data_col17[17] <= data_col17[16];

   data_col18[1] <= data[147];
   data_col18[2] <= data_col18[1];
   data_col18[3] <= data_col18[2];
   data_col18[4] <= data_col18[3];
   data_col18[5] <= data_col18[4];
   data_col18[6] <= data_col18[5];
   data_col18[7] <= data_col18[6];
   data_col18[8] <= data_col18[7];
   data_col18[9] <= data_col18[8];
   data_col18[10] <= data_col18[9];
   data_col18[11] <= data_col18[10];
   data_col18[12] <= data_col18[11];
   data_col18[13] <= data_col18[12];
   data_col18[14] <= data_col18[13];
   data_col18[15] <= data_col18[14];
   data_col18[16] <= data_col18[15];
   data_col18[17] <= data_col18[16];
   data_col18[18] <= data_col18[17];

   data_col19[1] <= data[146];
   data_col19[2] <= data_col19[1];
   data_col19[3] <= data_col19[2];
   data_col19[4] <= data_col19[3];
   data_col19[5] <= data_col19[4];
   data_col19[6] <= data_col19[5];
   data_col19[7] <= data_col19[6];
   data_col19[8] <= data_col19[7];
   data_col19[9] <= data_col19[8];
   data_col19[10] <= data_col19[9];
   data_col19[11] <= data_col19[10];
   data_col19[12] <= data_col19[11];
   data_col19[13] <= data_col19[12];
   data_col19[14] <= data_col19[13];
   data_col19[15] <= data_col19[14];
   data_col19[16] <= data_col19[15];
   data_col19[17] <= data_col19[16];
   data_col19[18] <= data_col19[17];
   data_col19[19] <= data_col19[18];

   data_col20[1] <= data[145];
   data_col20[2] <= data_col20[1];
   data_col20[3] <= data_col20[2];
   data_col20[4] <= data_col20[3];
   data_col20[5] <= data_col20[4];
   data_col20[6] <= data_col20[5];
   data_col20[7] <= data_col20[6];
   data_col20[8] <= data_col20[7];
   data_col20[9] <= data_col20[8];
   data_col20[10] <= data_col20[9];
   data_col20[11] <= data_col20[10];
   data_col20[12] <= data_col20[11];
   data_col20[13] <= data_col20[12];
   data_col20[14] <= data_col20[13];
   data_col20[15] <= data_col20[14];
   data_col20[16] <= data_col20[15];
   data_col20[17] <= data_col20[16];
   data_col20[18] <= data_col20[17];
   data_col20[19] <= data_col20[18];
   data_col20[20] <= data_col20[19];

   data_col21[1] <= data[144];
   data_col21[2] <= data_col21[1];
   data_col21[3] <= data_col21[2];
   data_col21[4] <= data_col21[3];
   data_col21[5] <= data_col21[4];
   data_col21[6] <= data_col21[5];
   data_col21[7] <= data_col21[6];
   data_col21[8] <= data_col21[7];
   data_col21[9] <= data_col21[8];
   data_col21[10] <= data_col21[9];
   data_col21[11] <= data_col21[10];
   data_col21[12] <= data_col21[11];
   data_col21[13] <= data_col21[12];
   data_col21[14] <= data_col21[13];
   data_col21[15] <= data_col21[14];
   data_col21[16] <= data_col21[15];
   data_col21[17] <= data_col21[16];
   data_col21[18] <= data_col21[17];
   data_col21[19] <= data_col21[18];
   data_col21[20] <= data_col21[19];
   data_col21[21] <= data_col21[20];

   data_col22[1] <= data[143];
   data_col22[2] <= data_col22[1];
   data_col22[3] <= data_col22[2];
   data_col22[4] <= data_col22[3];
   data_col22[5] <= data_col22[4];
   data_col22[6] <= data_col22[5];
   data_col22[7] <= data_col22[6];
   data_col22[8] <= data_col22[7];
   data_col22[9] <= data_col22[8];
   data_col22[10] <= data_col22[9];
   data_col22[11] <= data_col22[10];
   data_col22[12] <= data_col22[11];
   data_col22[13] <= data_col22[12];
   data_col22[14] <= data_col22[13];
   data_col22[15] <= data_col22[14];
   data_col22[16] <= data_col22[15];
   data_col22[17] <= data_col22[16];
   data_col22[18] <= data_col22[17];
   data_col22[19] <= data_col22[18];
   data_col22[20] <= data_col22[19];
   data_col22[21] <= data_col22[20];
   data_col22[22] <= data_col22[21];

   data_col23[1] <= data[142];
   data_col23[2] <= data_col23[1];
   data_col23[3] <= data_col23[2];
   data_col23[4] <= data_col23[3];
   data_col23[5] <= data_col23[4];
   data_col23[6] <= data_col23[5];
   data_col23[7] <= data_col23[6];
   data_col23[8] <= data_col23[7];
   data_col23[9] <= data_col23[8];
   data_col23[10] <= data_col23[9];
   data_col23[11] <= data_col23[10];
   data_col23[12] <= data_col23[11];
   data_col23[13] <= data_col23[12];
   data_col23[14] <= data_col23[13];
   data_col23[15] <= data_col23[14];
   data_col23[16] <= data_col23[15];
   data_col23[17] <= data_col23[16];
   data_col23[18] <= data_col23[17];
   data_col23[19] <= data_col23[18];
   data_col23[20] <= data_col23[19];
   data_col23[21] <= data_col23[20];
   data_col23[22] <= data_col23[21];
   data_col23[23] <= data_col23[22];

   data_col24[1] <= data[141];
   data_col24[2] <= data_col24[1];
   data_col24[3] <= data_col24[2];
   data_col24[4] <= data_col24[3];
   data_col24[5] <= data_col24[4];
   data_col24[6] <= data_col24[5];
   data_col24[7] <= data_col24[6];
   data_col24[8] <= data_col24[7];
   data_col24[9] <= data_col24[8];
   data_col24[10] <= data_col24[9];
   data_col24[11] <= data_col24[10];
   data_col24[12] <= data_col24[11];
   data_col24[13] <= data_col24[12];
   data_col24[14] <= data_col24[13];
   data_col24[15] <= data_col24[14];
   data_col24[16] <= data_col24[15];
   data_col24[17] <= data_col24[16];
   data_col24[18] <= data_col24[17];
   data_col24[19] <= data_col24[18];
   data_col24[20] <= data_col24[19];
   data_col24[21] <= data_col24[20];
   data_col24[22] <= data_col24[21];
   data_col24[23] <= data_col24[22];
   data_col24[24] <= data_col24[23];

   data_col25[1] <= data[140];
   data_col25[2] <= data_col25[1];
   data_col25[3] <= data_col25[2];
   data_col25[4] <= data_col25[3];
   data_col25[5] <= data_col25[4];
   data_col25[6] <= data_col25[5];
   data_col25[7] <= data_col25[6];
   data_col25[8] <= data_col25[7];
   data_col25[9] <= data_col25[8];
   data_col25[10] <= data_col25[9];
   data_col25[11] <= data_col25[10];
   data_col25[12] <= data_col25[11];
   data_col25[13] <= data_col25[12];
   data_col25[14] <= data_col25[13];
   data_col25[15] <= data_col25[14];
   data_col25[16] <= data_col25[15];
   data_col25[17] <= data_col25[16];
   data_col25[18] <= data_col25[17];
   data_col25[19] <= data_col25[18];
   data_col25[20] <= data_col25[19];
   data_col25[21] <= data_col25[20];
   data_col25[22] <= data_col25[21];
   data_col25[23] <= data_col25[22];
   data_col25[24] <= data_col25[23];
   data_col25[25] <= data_col25[24];

   data_col26[1] <= data[139];
   data_col26[2] <= data_col26[1];
   data_col26[3] <= data_col26[2];
   data_col26[4] <= data_col26[3];
   data_col26[5] <= data_col26[4];
   data_col26[6] <= data_col26[5];
   data_col26[7] <= data_col26[6];
   data_col26[8] <= data_col26[7];
   data_col26[9] <= data_col26[8];
   data_col26[10] <= data_col26[9];
   data_col26[11] <= data_col26[10];
   data_col26[12] <= data_col26[11];
   data_col26[13] <= data_col26[12];
   data_col26[14] <= data_col26[13];
   data_col26[15] <= data_col26[14];
   data_col26[16] <= data_col26[15];
   data_col26[17] <= data_col26[16];
   data_col26[18] <= data_col26[17];
   data_col26[19] <= data_col26[18];
   data_col26[20] <= data_col26[19];
   data_col26[21] <= data_col26[20];
   data_col26[22] <= data_col26[21];
   data_col26[23] <= data_col26[22];
   data_col26[24] <= data_col26[23];
   data_col26[25] <= data_col26[24];
   data_col26[26] <= data_col26[25];

   data_col27[1] <= data[138];
   data_col27[2] <= data_col27[1];
   data_col27[3] <= data_col27[2];
   data_col27[4] <= data_col27[3];
   data_col27[5] <= data_col27[4];
   data_col27[6] <= data_col27[5];
   data_col27[7] <= data_col27[6];
   data_col27[8] <= data_col27[7];
   data_col27[9] <= data_col27[8];
   data_col27[10] <= data_col27[9];
   data_col27[11] <= data_col27[10];
   data_col27[12] <= data_col27[11];
   data_col27[13] <= data_col27[12];
   data_col27[14] <= data_col27[13];
   data_col27[15] <= data_col27[14];
   data_col27[16] <= data_col27[15];
   data_col27[17] <= data_col27[16];
   data_col27[18] <= data_col27[17];
   data_col27[19] <= data_col27[18];
   data_col27[20] <= data_col27[19];
   data_col27[21] <= data_col27[20];
   data_col27[22] <= data_col27[21];
   data_col27[23] <= data_col27[22];
   data_col27[24] <= data_col27[23];
   data_col27[25] <= data_col27[24];
   data_col27[26] <= data_col27[25];
   data_col27[27] <= data_col27[26];

   data_col28[1] <= data[137];
   data_col28[2] <= data_col28[1];
   data_col28[3] <= data_col28[2];
   data_col28[4] <= data_col28[3];
   data_col28[5] <= data_col28[4];
   data_col28[6] <= data_col28[5];
   data_col28[7] <= data_col28[6];
   data_col28[8] <= data_col28[7];
   data_col28[9] <= data_col28[8];
   data_col28[10] <= data_col28[9];
   data_col28[11] <= data_col28[10];
   data_col28[12] <= data_col28[11];
   data_col28[13] <= data_col28[12];
   data_col28[14] <= data_col28[13];
   data_col28[15] <= data_col28[14];
   data_col28[16] <= data_col28[15];
   data_col28[17] <= data_col28[16];
   data_col28[18] <= data_col28[17];
   data_col28[19] <= data_col28[18];
   data_col28[20] <= data_col28[19];
   data_col28[21] <= data_col28[20];
   data_col28[22] <= data_col28[21];
   data_col28[23] <= data_col28[22];
   data_col28[24] <= data_col28[23];
   data_col28[25] <= data_col28[24];
   data_col28[26] <= data_col28[25];
   data_col28[27] <= data_col28[26];
   data_col28[28] <= data_col28[27];

   data_col29[1] <= data[136];
   data_col29[2] <= data_col29[1];
   data_col29[3] <= data_col29[2];
   data_col29[4] <= data_col29[3];
   data_col29[5] <= data_col29[4];
   data_col29[6] <= data_col29[5];
   data_col29[7] <= data_col29[6];
   data_col29[8] <= data_col29[7];
   data_col29[9] <= data_col29[8];
   data_col29[10] <= data_col29[9];
   data_col29[11] <= data_col29[10];
   data_col29[12] <= data_col29[11];
   data_col29[13] <= data_col29[12];
   data_col29[14] <= data_col29[13];
   data_col29[15] <= data_col29[14];
   data_col29[16] <= data_col29[15];
   data_col29[17] <= data_col29[16];
   data_col29[18] <= data_col29[17];
   data_col29[19] <= data_col29[18];
   data_col29[20] <= data_col29[19];
   data_col29[21] <= data_col29[20];
   data_col29[22] <= data_col29[21];
   data_col29[23] <= data_col29[22];
   data_col29[24] <= data_col29[23];
   data_col29[25] <= data_col29[24];
   data_col29[26] <= data_col29[25];
   data_col29[27] <= data_col29[26];
   data_col29[28] <= data_col29[27];
   data_col29[29] <= data_col29[28];

   data_col30[1] <= data[135];
   data_col30[2] <= data_col30[1];
   data_col30[3] <= data_col30[2];
   data_col30[4] <= data_col30[3];
   data_col30[5] <= data_col30[4];
   data_col30[6] <= data_col30[5];
   data_col30[7] <= data_col30[6];
   data_col30[8] <= data_col30[7];
   data_col30[9] <= data_col30[8];
   data_col30[10] <= data_col30[9];
   data_col30[11] <= data_col30[10];
   data_col30[12] <= data_col30[11];
   data_col30[13] <= data_col30[12];
   data_col30[14] <= data_col30[13];
   data_col30[15] <= data_col30[14];
   data_col30[16] <= data_col30[15];
   data_col30[17] <= data_col30[16];
   data_col30[18] <= data_col30[17];
   data_col30[19] <= data_col30[18];
   data_col30[20] <= data_col30[19];
   data_col30[21] <= data_col30[20];
   data_col30[22] <= data_col30[21];
   data_col30[23] <= data_col30[22];
   data_col30[24] <= data_col30[23];
   data_col30[25] <= data_col30[24];
   data_col30[26] <= data_col30[25];
   data_col30[27] <= data_col30[26];
   data_col30[28] <= data_col30[27];
   data_col30[29] <= data_col30[28];
   data_col30[30] <= data_col30[29];

   data_col31[1] <= data[134];
   data_col31[2] <= data_col31[1];
   data_col31[3] <= data_col31[2];
   data_col31[4] <= data_col31[3];
   data_col31[5] <= data_col31[4];
   data_col31[6] <= data_col31[5];
   data_col31[7] <= data_col31[6];
   data_col31[8] <= data_col31[7];
   data_col31[9] <= data_col31[8];
   data_col31[10] <= data_col31[9];
   data_col31[11] <= data_col31[10];
   data_col31[12] <= data_col31[11];
   data_col31[13] <= data_col31[12];
   data_col31[14] <= data_col31[13];
   data_col31[15] <= data_col31[14];
   data_col31[16] <= data_col31[15];
   data_col31[17] <= data_col31[16];
   data_col31[18] <= data_col31[17];
   data_col31[19] <= data_col31[18];
   data_col31[20] <= data_col31[19];
   data_col31[21] <= data_col31[20];
   data_col31[22] <= data_col31[21];
   data_col31[23] <= data_col31[22];
   data_col31[24] <= data_col31[23];
   data_col31[25] <= data_col31[24];
   data_col31[26] <= data_col31[25];
   data_col31[27] <= data_col31[26];
   data_col31[28] <= data_col31[27];
   data_col31[29] <= data_col31[28];
   data_col31[30] <= data_col31[29];
   data_col31[31] <= data_col31[30];

   data_col32[1] <= data[133];
   data_col32[2] <= data_col32[1];
   data_col32[3] <= data_col32[2];
   data_col32[4] <= data_col32[3];
   data_col32[5] <= data_col32[4];
   data_col32[6] <= data_col32[5];
   data_col32[7] <= data_col32[6];
   data_col32[8] <= data_col32[7];
   data_col32[9] <= data_col32[8];
   data_col32[10] <= data_col32[9];
   data_col32[11] <= data_col32[10];
   data_col32[12] <= data_col32[11];
   data_col32[13] <= data_col32[12];
   data_col32[14] <= data_col32[13];
   data_col32[15] <= data_col32[14];
   data_col32[16] <= data_col32[15];
   data_col32[17] <= data_col32[16];
   data_col32[18] <= data_col32[17];
   data_col32[19] <= data_col32[18];
   data_col32[20] <= data_col32[19];
   data_col32[21] <= data_col32[20];
   data_col32[22] <= data_col32[21];
   data_col32[23] <= data_col32[22];
   data_col32[24] <= data_col32[23];
   data_col32[25] <= data_col32[24];
   data_col32[26] <= data_col32[25];
   data_col32[27] <= data_col32[26];
   data_col32[28] <= data_col32[27];
   data_col32[29] <= data_col32[28];
   data_col32[30] <= data_col32[29];
   data_col32[31] <= data_col32[30];
   data_col32[32] <= data_col32[31];

   data_col33[1] <= data[132];
   data_col33[2] <= data_col33[1];
   data_col33[3] <= data_col33[2];
   data_col33[4] <= data_col33[3];
   data_col33[5] <= data_col33[4];
   data_col33[6] <= data_col33[5];
   data_col33[7] <= data_col33[6];
   data_col33[8] <= data_col33[7];
   data_col33[9] <= data_col33[8];
   data_col33[10] <= data_col33[9];
   data_col33[11] <= data_col33[10];
   data_col33[12] <= data_col33[11];
   data_col33[13] <= data_col33[12];
   data_col33[14] <= data_col33[13];
   data_col33[15] <= data_col33[14];
   data_col33[16] <= data_col33[15];
   data_col33[17] <= data_col33[16];
   data_col33[18] <= data_col33[17];
   data_col33[19] <= data_col33[18];
   data_col33[20] <= data_col33[19];
   data_col33[21] <= data_col33[20];
   data_col33[22] <= data_col33[21];
   data_col33[23] <= data_col33[22];
   data_col33[24] <= data_col33[23];
   data_col33[25] <= data_col33[24];
   data_col33[26] <= data_col33[25];
   data_col33[27] <= data_col33[26];
   data_col33[28] <= data_col33[27];
   data_col33[29] <= data_col33[28];
   data_col33[30] <= data_col33[29];
   data_col33[31] <= data_col33[30];
   data_col33[32] <= data_col33[31];
   data_col33[33] <= data_col33[32];

   data_col34[1] <= data[131];
   data_col34[2] <= data_col34[1];
   data_col34[3] <= data_col34[2];
   data_col34[4] <= data_col34[3];
   data_col34[5] <= data_col34[4];
   data_col34[6] <= data_col34[5];
   data_col34[7] <= data_col34[6];
   data_col34[8] <= data_col34[7];
   data_col34[9] <= data_col34[8];
   data_col34[10] <= data_col34[9];
   data_col34[11] <= data_col34[10];
   data_col34[12] <= data_col34[11];
   data_col34[13] <= data_col34[12];
   data_col34[14] <= data_col34[13];
   data_col34[15] <= data_col34[14];
   data_col34[16] <= data_col34[15];
   data_col34[17] <= data_col34[16];
   data_col34[18] <= data_col34[17];
   data_col34[19] <= data_col34[18];
   data_col34[20] <= data_col34[19];
   data_col34[21] <= data_col34[20];
   data_col34[22] <= data_col34[21];
   data_col34[23] <= data_col34[22];
   data_col34[24] <= data_col34[23];
   data_col34[25] <= data_col34[24];
   data_col34[26] <= data_col34[25];
   data_col34[27] <= data_col34[26];
   data_col34[28] <= data_col34[27];
   data_col34[29] <= data_col34[28];
   data_col34[30] <= data_col34[29];
   data_col34[31] <= data_col34[30];
   data_col34[32] <= data_col34[31];
   data_col34[33] <= data_col34[32];
   data_col34[34] <= data_col34[33];

   data_col35[1] <= data[130];
   data_col35[2] <= data_col35[1];
   data_col35[3] <= data_col35[2];
   data_col35[4] <= data_col35[3];
   data_col35[5] <= data_col35[4];
   data_col35[6] <= data_col35[5];
   data_col35[7] <= data_col35[6];
   data_col35[8] <= data_col35[7];
   data_col35[9] <= data_col35[8];
   data_col35[10] <= data_col35[9];
   data_col35[11] <= data_col35[10];
   data_col35[12] <= data_col35[11];
   data_col35[13] <= data_col35[12];
   data_col35[14] <= data_col35[13];
   data_col35[15] <= data_col35[14];
   data_col35[16] <= data_col35[15];
   data_col35[17] <= data_col35[16];
   data_col35[18] <= data_col35[17];
   data_col35[19] <= data_col35[18];
   data_col35[20] <= data_col35[19];
   data_col35[21] <= data_col35[20];
   data_col35[22] <= data_col35[21];
   data_col35[23] <= data_col35[22];
   data_col35[24] <= data_col35[23];
   data_col35[25] <= data_col35[24];
   data_col35[26] <= data_col35[25];
   data_col35[27] <= data_col35[26];
   data_col35[28] <= data_col35[27];
   data_col35[29] <= data_col35[28];
   data_col35[30] <= data_col35[29];
   data_col35[31] <= data_col35[30];
   data_col35[32] <= data_col35[31];
   data_col35[33] <= data_col35[32];
   data_col35[34] <= data_col35[33];
   data_col35[35] <= data_col35[34];

   data_col36[1] <= data[129];
   data_col36[2] <= data_col36[1];
   data_col36[3] <= data_col36[2];
   data_col36[4] <= data_col36[3];
   data_col36[5] <= data_col36[4];
   data_col36[6] <= data_col36[5];
   data_col36[7] <= data_col36[6];
   data_col36[8] <= data_col36[7];
   data_col36[9] <= data_col36[8];
   data_col36[10] <= data_col36[9];
   data_col36[11] <= data_col36[10];
   data_col36[12] <= data_col36[11];
   data_col36[13] <= data_col36[12];
   data_col36[14] <= data_col36[13];
   data_col36[15] <= data_col36[14];
   data_col36[16] <= data_col36[15];
   data_col36[17] <= data_col36[16];
   data_col36[18] <= data_col36[17];
   data_col36[19] <= data_col36[18];
   data_col36[20] <= data_col36[19];
   data_col36[21] <= data_col36[20];
   data_col36[22] <= data_col36[21];
   data_col36[23] <= data_col36[22];
   data_col36[24] <= data_col36[23];
   data_col36[25] <= data_col36[24];
   data_col36[26] <= data_col36[25];
   data_col36[27] <= data_col36[26];
   data_col36[28] <= data_col36[27];
   data_col36[29] <= data_col36[28];
   data_col36[30] <= data_col36[29];
   data_col36[31] <= data_col36[30];
   data_col36[32] <= data_col36[31];
   data_col36[33] <= data_col36[32];
   data_col36[34] <= data_col36[33];
   data_col36[35] <= data_col36[34];
   data_col36[36] <= data_col36[35];

   data_col37[1] <= data[128];
   data_col37[2] <= data_col37[1];
   data_col37[3] <= data_col37[2];
   data_col37[4] <= data_col37[3];
   data_col37[5] <= data_col37[4];
   data_col37[6] <= data_col37[5];
   data_col37[7] <= data_col37[6];
   data_col37[8] <= data_col37[7];
   data_col37[9] <= data_col37[8];
   data_col37[10] <= data_col37[9];
   data_col37[11] <= data_col37[10];
   data_col37[12] <= data_col37[11];
   data_col37[13] <= data_col37[12];
   data_col37[14] <= data_col37[13];
   data_col37[15] <= data_col37[14];
   data_col37[16] <= data_col37[15];
   data_col37[17] <= data_col37[16];
   data_col37[18] <= data_col37[17];
   data_col37[19] <= data_col37[18];
   data_col37[20] <= data_col37[19];
   data_col37[21] <= data_col37[20];
   data_col37[22] <= data_col37[21];
   data_col37[23] <= data_col37[22];
   data_col37[24] <= data_col37[23];
   data_col37[25] <= data_col37[24];
   data_col37[26] <= data_col37[25];
   data_col37[27] <= data_col37[26];
   data_col37[28] <= data_col37[27];
   data_col37[29] <= data_col37[28];
   data_col37[30] <= data_col37[29];
   data_col37[31] <= data_col37[30];
   data_col37[32] <= data_col37[31];
   data_col37[33] <= data_col37[32];
   data_col37[34] <= data_col37[33];
   data_col37[35] <= data_col37[34];
   data_col37[36] <= data_col37[35];
   data_col37[37] <= data_col37[36];

   data_col38[1] <= data[127];
   data_col38[2] <= data_col38[1];
   data_col38[3] <= data_col38[2];
   data_col38[4] <= data_col38[3];
   data_col38[5] <= data_col38[4];
   data_col38[6] <= data_col38[5];
   data_col38[7] <= data_col38[6];
   data_col38[8] <= data_col38[7];
   data_col38[9] <= data_col38[8];
   data_col38[10] <= data_col38[9];
   data_col38[11] <= data_col38[10];
   data_col38[12] <= data_col38[11];
   data_col38[13] <= data_col38[12];
   data_col38[14] <= data_col38[13];
   data_col38[15] <= data_col38[14];
   data_col38[16] <= data_col38[15];
   data_col38[17] <= data_col38[16];
   data_col38[18] <= data_col38[17];
   data_col38[19] <= data_col38[18];
   data_col38[20] <= data_col38[19];
   data_col38[21] <= data_col38[20];
   data_col38[22] <= data_col38[21];
   data_col38[23] <= data_col38[22];
   data_col38[24] <= data_col38[23];
   data_col38[25] <= data_col38[24];
   data_col38[26] <= data_col38[25];
   data_col38[27] <= data_col38[26];
   data_col38[28] <= data_col38[27];
   data_col38[29] <= data_col38[28];
   data_col38[30] <= data_col38[29];
   data_col38[31] <= data_col38[30];
   data_col38[32] <= data_col38[31];
   data_col38[33] <= data_col38[32];
   data_col38[34] <= data_col38[33];
   data_col38[35] <= data_col38[34];
   data_col38[36] <= data_col38[35];
   data_col38[37] <= data_col38[36];
   data_col38[38] <= data_col38[37];

   data_col39[1] <= data[126];
   data_col39[2] <= data_col39[1];
   data_col39[3] <= data_col39[2];
   data_col39[4] <= data_col39[3];
   data_col39[5] <= data_col39[4];
   data_col39[6] <= data_col39[5];
   data_col39[7] <= data_col39[6];
   data_col39[8] <= data_col39[7];
   data_col39[9] <= data_col39[8];
   data_col39[10] <= data_col39[9];
   data_col39[11] <= data_col39[10];
   data_col39[12] <= data_col39[11];
   data_col39[13] <= data_col39[12];
   data_col39[14] <= data_col39[13];
   data_col39[15] <= data_col39[14];
   data_col39[16] <= data_col39[15];
   data_col39[17] <= data_col39[16];
   data_col39[18] <= data_col39[17];
   data_col39[19] <= data_col39[18];
   data_col39[20] <= data_col39[19];
   data_col39[21] <= data_col39[20];
   data_col39[22] <= data_col39[21];
   data_col39[23] <= data_col39[22];
   data_col39[24] <= data_col39[23];
   data_col39[25] <= data_col39[24];
   data_col39[26] <= data_col39[25];
   data_col39[27] <= data_col39[26];
   data_col39[28] <= data_col39[27];
   data_col39[29] <= data_col39[28];
   data_col39[30] <= data_col39[29];
   data_col39[31] <= data_col39[30];
   data_col39[32] <= data_col39[31];
   data_col39[33] <= data_col39[32];
   data_col39[34] <= data_col39[33];
   data_col39[35] <= data_col39[34];
   data_col39[36] <= data_col39[35];
   data_col39[37] <= data_col39[36];
   data_col39[38] <= data_col39[37];
   data_col39[39] <= data_col39[38];

   data_col40[1] <= data[125];
   data_col40[2] <= data_col40[1];
   data_col40[3] <= data_col40[2];
   data_col40[4] <= data_col40[3];
   data_col40[5] <= data_col40[4];
   data_col40[6] <= data_col40[5];
   data_col40[7] <= data_col40[6];
   data_col40[8] <= data_col40[7];
   data_col40[9] <= data_col40[8];
   data_col40[10] <= data_col40[9];
   data_col40[11] <= data_col40[10];
   data_col40[12] <= data_col40[11];
   data_col40[13] <= data_col40[12];
   data_col40[14] <= data_col40[13];
   data_col40[15] <= data_col40[14];
   data_col40[16] <= data_col40[15];
   data_col40[17] <= data_col40[16];
   data_col40[18] <= data_col40[17];
   data_col40[19] <= data_col40[18];
   data_col40[20] <= data_col40[19];
   data_col40[21] <= data_col40[20];
   data_col40[22] <= data_col40[21];
   data_col40[23] <= data_col40[22];
   data_col40[24] <= data_col40[23];
   data_col40[25] <= data_col40[24];
   data_col40[26] <= data_col40[25];
   data_col40[27] <= data_col40[26];
   data_col40[28] <= data_col40[27];
   data_col40[29] <= data_col40[28];
   data_col40[30] <= data_col40[29];
   data_col40[31] <= data_col40[30];
   data_col40[32] <= data_col40[31];
   data_col40[33] <= data_col40[32];
   data_col40[34] <= data_col40[33];
   data_col40[35] <= data_col40[34];
   data_col40[36] <= data_col40[35];
   data_col40[37] <= data_col40[36];
   data_col40[38] <= data_col40[37];
   data_col40[39] <= data_col40[38];
   data_col40[40] <= data_col40[39];

   data_col41[1] <= data[124];
   data_col41[2] <= data_col41[1];
   data_col41[3] <= data_col41[2];
   data_col41[4] <= data_col41[3];
   data_col41[5] <= data_col41[4];
   data_col41[6] <= data_col41[5];
   data_col41[7] <= data_col41[6];
   data_col41[8] <= data_col41[7];
   data_col41[9] <= data_col41[8];
   data_col41[10] <= data_col41[9];
   data_col41[11] <= data_col41[10];
   data_col41[12] <= data_col41[11];
   data_col41[13] <= data_col41[12];
   data_col41[14] <= data_col41[13];
   data_col41[15] <= data_col41[14];
   data_col41[16] <= data_col41[15];
   data_col41[17] <= data_col41[16];
   data_col41[18] <= data_col41[17];
   data_col41[19] <= data_col41[18];
   data_col41[20] <= data_col41[19];
   data_col41[21] <= data_col41[20];
   data_col41[22] <= data_col41[21];
   data_col41[23] <= data_col41[22];
   data_col41[24] <= data_col41[23];
   data_col41[25] <= data_col41[24];
   data_col41[26] <= data_col41[25];
   data_col41[27] <= data_col41[26];
   data_col41[28] <= data_col41[27];
   data_col41[29] <= data_col41[28];
   data_col41[30] <= data_col41[29];
   data_col41[31] <= data_col41[30];
   data_col41[32] <= data_col41[31];
   data_col41[33] <= data_col41[32];
   data_col41[34] <= data_col41[33];
   data_col41[35] <= data_col41[34];
   data_col41[36] <= data_col41[35];
   data_col41[37] <= data_col41[36];
   data_col41[38] <= data_col41[37];
   data_col41[39] <= data_col41[38];
   data_col41[40] <= data_col41[39];
   data_col41[41] <= data_col41[40];

   data_col42[1] <= data[123];
   data_col42[2] <= data_col42[1];
   data_col42[3] <= data_col42[2];
   data_col42[4] <= data_col42[3];
   data_col42[5] <= data_col42[4];
   data_col42[6] <= data_col42[5];
   data_col42[7] <= data_col42[6];
   data_col42[8] <= data_col42[7];
   data_col42[9] <= data_col42[8];
   data_col42[10] <= data_col42[9];
   data_col42[11] <= data_col42[10];
   data_col42[12] <= data_col42[11];
   data_col42[13] <= data_col42[12];
   data_col42[14] <= data_col42[13];
   data_col42[15] <= data_col42[14];
   data_col42[16] <= data_col42[15];
   data_col42[17] <= data_col42[16];
   data_col42[18] <= data_col42[17];
   data_col42[19] <= data_col42[18];
   data_col42[20] <= data_col42[19];
   data_col42[21] <= data_col42[20];
   data_col42[22] <= data_col42[21];
   data_col42[23] <= data_col42[22];
   data_col42[24] <= data_col42[23];
   data_col42[25] <= data_col42[24];
   data_col42[26] <= data_col42[25];
   data_col42[27] <= data_col42[26];
   data_col42[28] <= data_col42[27];
   data_col42[29] <= data_col42[28];
   data_col42[30] <= data_col42[29];
   data_col42[31] <= data_col42[30];
   data_col42[32] <= data_col42[31];
   data_col42[33] <= data_col42[32];
   data_col42[34] <= data_col42[33];
   data_col42[35] <= data_col42[34];
   data_col42[36] <= data_col42[35];
   data_col42[37] <= data_col42[36];
   data_col42[38] <= data_col42[37];
   data_col42[39] <= data_col42[38];
   data_col42[40] <= data_col42[39];
   data_col42[41] <= data_col42[40];
   data_col42[42] <= data_col42[41];

   data_col43[1] <= data[122];
   data_col43[2] <= data_col43[1];
   data_col43[3] <= data_col43[2];
   data_col43[4] <= data_col43[3];
   data_col43[5] <= data_col43[4];
   data_col43[6] <= data_col43[5];
   data_col43[7] <= data_col43[6];
   data_col43[8] <= data_col43[7];
   data_col43[9] <= data_col43[8];
   data_col43[10] <= data_col43[9];
   data_col43[11] <= data_col43[10];
   data_col43[12] <= data_col43[11];
   data_col43[13] <= data_col43[12];
   data_col43[14] <= data_col43[13];
   data_col43[15] <= data_col43[14];
   data_col43[16] <= data_col43[15];
   data_col43[17] <= data_col43[16];
   data_col43[18] <= data_col43[17];
   data_col43[19] <= data_col43[18];
   data_col43[20] <= data_col43[19];
   data_col43[21] <= data_col43[20];
   data_col43[22] <= data_col43[21];
   data_col43[23] <= data_col43[22];
   data_col43[24] <= data_col43[23];
   data_col43[25] <= data_col43[24];
   data_col43[26] <= data_col43[25];
   data_col43[27] <= data_col43[26];
   data_col43[28] <= data_col43[27];
   data_col43[29] <= data_col43[28];
   data_col43[30] <= data_col43[29];
   data_col43[31] <= data_col43[30];
   data_col43[32] <= data_col43[31];
   data_col43[33] <= data_col43[32];
   data_col43[34] <= data_col43[33];
   data_col43[35] <= data_col43[34];
   data_col43[36] <= data_col43[35];
   data_col43[37] <= data_col43[36];
   data_col43[38] <= data_col43[37];
   data_col43[39] <= data_col43[38];
   data_col43[40] <= data_col43[39];
   data_col43[41] <= data_col43[40];
   data_col43[42] <= data_col43[41];
   data_col43[43] <= data_col43[42];

   data_col44[1] <= data[121];
   data_col44[2] <= data_col44[1];
   data_col44[3] <= data_col44[2];
   data_col44[4] <= data_col44[3];
   data_col44[5] <= data_col44[4];
   data_col44[6] <= data_col44[5];
   data_col44[7] <= data_col44[6];
   data_col44[8] <= data_col44[7];
   data_col44[9] <= data_col44[8];
   data_col44[10] <= data_col44[9];
   data_col44[11] <= data_col44[10];
   data_col44[12] <= data_col44[11];
   data_col44[13] <= data_col44[12];
   data_col44[14] <= data_col44[13];
   data_col44[15] <= data_col44[14];
   data_col44[16] <= data_col44[15];
   data_col44[17] <= data_col44[16];
   data_col44[18] <= data_col44[17];
   data_col44[19] <= data_col44[18];
   data_col44[20] <= data_col44[19];
   data_col44[21] <= data_col44[20];
   data_col44[22] <= data_col44[21];
   data_col44[23] <= data_col44[22];
   data_col44[24] <= data_col44[23];
   data_col44[25] <= data_col44[24];
   data_col44[26] <= data_col44[25];
   data_col44[27] <= data_col44[26];
   data_col44[28] <= data_col44[27];
   data_col44[29] <= data_col44[28];
   data_col44[30] <= data_col44[29];
   data_col44[31] <= data_col44[30];
   data_col44[32] <= data_col44[31];
   data_col44[33] <= data_col44[32];
   data_col44[34] <= data_col44[33];
   data_col44[35] <= data_col44[34];
   data_col44[36] <= data_col44[35];
   data_col44[37] <= data_col44[36];
   data_col44[38] <= data_col44[37];
   data_col44[39] <= data_col44[38];
   data_col44[40] <= data_col44[39];
   data_col44[41] <= data_col44[40];
   data_col44[42] <= data_col44[41];
   data_col44[43] <= data_col44[42];
   data_col44[44] <= data_col44[43];

   data_col45[1] <= data[120];
   data_col45[2] <= data_col45[1];
   data_col45[3] <= data_col45[2];
   data_col45[4] <= data_col45[3];
   data_col45[5] <= data_col45[4];
   data_col45[6] <= data_col45[5];
   data_col45[7] <= data_col45[6];
   data_col45[8] <= data_col45[7];
   data_col45[9] <= data_col45[8];
   data_col45[10] <= data_col45[9];
   data_col45[11] <= data_col45[10];
   data_col45[12] <= data_col45[11];
   data_col45[13] <= data_col45[12];
   data_col45[14] <= data_col45[13];
   data_col45[15] <= data_col45[14];
   data_col45[16] <= data_col45[15];
   data_col45[17] <= data_col45[16];
   data_col45[18] <= data_col45[17];
   data_col45[19] <= data_col45[18];
   data_col45[20] <= data_col45[19];
   data_col45[21] <= data_col45[20];
   data_col45[22] <= data_col45[21];
   data_col45[23] <= data_col45[22];
   data_col45[24] <= data_col45[23];
   data_col45[25] <= data_col45[24];
   data_col45[26] <= data_col45[25];
   data_col45[27] <= data_col45[26];
   data_col45[28] <= data_col45[27];
   data_col45[29] <= data_col45[28];
   data_col45[30] <= data_col45[29];
   data_col45[31] <= data_col45[30];
   data_col45[32] <= data_col45[31];
   data_col45[33] <= data_col45[32];
   data_col45[34] <= data_col45[33];
   data_col45[35] <= data_col45[34];
   data_col45[36] <= data_col45[35];
   data_col45[37] <= data_col45[36];
   data_col45[38] <= data_col45[37];
   data_col45[39] <= data_col45[38];
   data_col45[40] <= data_col45[39];
   data_col45[41] <= data_col45[40];
   data_col45[42] <= data_col45[41];
   data_col45[43] <= data_col45[42];
   data_col45[44] <= data_col45[43];
   data_col45[45] <= data_col45[44];

   data_col46[1] <= data[119];
   data_col46[2] <= data_col46[1];
   data_col46[3] <= data_col46[2];
   data_col46[4] <= data_col46[3];
   data_col46[5] <= data_col46[4];
   data_col46[6] <= data_col46[5];
   data_col46[7] <= data_col46[6];
   data_col46[8] <= data_col46[7];
   data_col46[9] <= data_col46[8];
   data_col46[10] <= data_col46[9];
   data_col46[11] <= data_col46[10];
   data_col46[12] <= data_col46[11];
   data_col46[13] <= data_col46[12];
   data_col46[14] <= data_col46[13];
   data_col46[15] <= data_col46[14];
   data_col46[16] <= data_col46[15];
   data_col46[17] <= data_col46[16];
   data_col46[18] <= data_col46[17];
   data_col46[19] <= data_col46[18];
   data_col46[20] <= data_col46[19];
   data_col46[21] <= data_col46[20];
   data_col46[22] <= data_col46[21];
   data_col46[23] <= data_col46[22];
   data_col46[24] <= data_col46[23];
   data_col46[25] <= data_col46[24];
   data_col46[26] <= data_col46[25];
   data_col46[27] <= data_col46[26];
   data_col46[28] <= data_col46[27];
   data_col46[29] <= data_col46[28];
   data_col46[30] <= data_col46[29];
   data_col46[31] <= data_col46[30];
   data_col46[32] <= data_col46[31];
   data_col46[33] <= data_col46[32];
   data_col46[34] <= data_col46[33];
   data_col46[35] <= data_col46[34];
   data_col46[36] <= data_col46[35];
   data_col46[37] <= data_col46[36];
   data_col46[38] <= data_col46[37];
   data_col46[39] <= data_col46[38];
   data_col46[40] <= data_col46[39];
   data_col46[41] <= data_col46[40];
   data_col46[42] <= data_col46[41];
   data_col46[43] <= data_col46[42];
   data_col46[44] <= data_col46[43];
   data_col46[45] <= data_col46[44];
   data_col46[46] <= data_col46[45];

   data_col47[1] <= data[118];
   data_col47[2] <= data_col47[1];
   data_col47[3] <= data_col47[2];
   data_col47[4] <= data_col47[3];
   data_col47[5] <= data_col47[4];
   data_col47[6] <= data_col47[5];
   data_col47[7] <= data_col47[6];
   data_col47[8] <= data_col47[7];
   data_col47[9] <= data_col47[8];
   data_col47[10] <= data_col47[9];
   data_col47[11] <= data_col47[10];
   data_col47[12] <= data_col47[11];
   data_col47[13] <= data_col47[12];
   data_col47[14] <= data_col47[13];
   data_col47[15] <= data_col47[14];
   data_col47[16] <= data_col47[15];
   data_col47[17] <= data_col47[16];
   data_col47[18] <= data_col47[17];
   data_col47[19] <= data_col47[18];
   data_col47[20] <= data_col47[19];
   data_col47[21] <= data_col47[20];
   data_col47[22] <= data_col47[21];
   data_col47[23] <= data_col47[22];
   data_col47[24] <= data_col47[23];
   data_col47[25] <= data_col47[24];
   data_col47[26] <= data_col47[25];
   data_col47[27] <= data_col47[26];
   data_col47[28] <= data_col47[27];
   data_col47[29] <= data_col47[28];
   data_col47[30] <= data_col47[29];
   data_col47[31] <= data_col47[30];
   data_col47[32] <= data_col47[31];
   data_col47[33] <= data_col47[32];
   data_col47[34] <= data_col47[33];
   data_col47[35] <= data_col47[34];
   data_col47[36] <= data_col47[35];
   data_col47[37] <= data_col47[36];
   data_col47[38] <= data_col47[37];
   data_col47[39] <= data_col47[38];
   data_col47[40] <= data_col47[39];
   data_col47[41] <= data_col47[40];
   data_col47[42] <= data_col47[41];
   data_col47[43] <= data_col47[42];
   data_col47[44] <= data_col47[43];
   data_col47[45] <= data_col47[44];
   data_col47[46] <= data_col47[45];
   data_col47[47] <= data_col47[46];

   data_col48[1] <= data[117];
   data_col48[2] <= data_col48[1];
   data_col48[3] <= data_col48[2];
   data_col48[4] <= data_col48[3];
   data_col48[5] <= data_col48[4];
   data_col48[6] <= data_col48[5];
   data_col48[7] <= data_col48[6];
   data_col48[8] <= data_col48[7];
   data_col48[9] <= data_col48[8];
   data_col48[10] <= data_col48[9];
   data_col48[11] <= data_col48[10];
   data_col48[12] <= data_col48[11];
   data_col48[13] <= data_col48[12];
   data_col48[14] <= data_col48[13];
   data_col48[15] <= data_col48[14];
   data_col48[16] <= data_col48[15];
   data_col48[17] <= data_col48[16];
   data_col48[18] <= data_col48[17];
   data_col48[19] <= data_col48[18];
   data_col48[20] <= data_col48[19];
   data_col48[21] <= data_col48[20];
   data_col48[22] <= data_col48[21];
   data_col48[23] <= data_col48[22];
   data_col48[24] <= data_col48[23];
   data_col48[25] <= data_col48[24];
   data_col48[26] <= data_col48[25];
   data_col48[27] <= data_col48[26];
   data_col48[28] <= data_col48[27];
   data_col48[29] <= data_col48[28];
   data_col48[30] <= data_col48[29];
   data_col48[31] <= data_col48[30];
   data_col48[32] <= data_col48[31];
   data_col48[33] <= data_col48[32];
   data_col48[34] <= data_col48[33];
   data_col48[35] <= data_col48[34];
   data_col48[36] <= data_col48[35];
   data_col48[37] <= data_col48[36];
   data_col48[38] <= data_col48[37];
   data_col48[39] <= data_col48[38];
   data_col48[40] <= data_col48[39];
   data_col48[41] <= data_col48[40];
   data_col48[42] <= data_col48[41];
   data_col48[43] <= data_col48[42];
   data_col48[44] <= data_col48[43];
   data_col48[45] <= data_col48[44];
   data_col48[46] <= data_col48[45];
   data_col48[47] <= data_col48[46];
   data_col48[48] <= data_col48[47];

   data_col49[1] <= data[116];
   data_col49[2] <= data_col49[1];
   data_col49[3] <= data_col49[2];
   data_col49[4] <= data_col49[3];
   data_col49[5] <= data_col49[4];
   data_col49[6] <= data_col49[5];
   data_col49[7] <= data_col49[6];
   data_col49[8] <= data_col49[7];
   data_col49[9] <= data_col49[8];
   data_col49[10] <= data_col49[9];
   data_col49[11] <= data_col49[10];
   data_col49[12] <= data_col49[11];
   data_col49[13] <= data_col49[12];
   data_col49[14] <= data_col49[13];
   data_col49[15] <= data_col49[14];
   data_col49[16] <= data_col49[15];
   data_col49[17] <= data_col49[16];
   data_col49[18] <= data_col49[17];
   data_col49[19] <= data_col49[18];
   data_col49[20] <= data_col49[19];
   data_col49[21] <= data_col49[20];
   data_col49[22] <= data_col49[21];
   data_col49[23] <= data_col49[22];
   data_col49[24] <= data_col49[23];
   data_col49[25] <= data_col49[24];
   data_col49[26] <= data_col49[25];
   data_col49[27] <= data_col49[26];
   data_col49[28] <= data_col49[27];
   data_col49[29] <= data_col49[28];
   data_col49[30] <= data_col49[29];
   data_col49[31] <= data_col49[30];
   data_col49[32] <= data_col49[31];
   data_col49[33] <= data_col49[32];
   data_col49[34] <= data_col49[33];
   data_col49[35] <= data_col49[34];
   data_col49[36] <= data_col49[35];
   data_col49[37] <= data_col49[36];
   data_col49[38] <= data_col49[37];
   data_col49[39] <= data_col49[38];
   data_col49[40] <= data_col49[39];
   data_col49[41] <= data_col49[40];
   data_col49[42] <= data_col49[41];
   data_col49[43] <= data_col49[42];
   data_col49[44] <= data_col49[43];
   data_col49[45] <= data_col49[44];
   data_col49[46] <= data_col49[45];
   data_col49[47] <= data_col49[46];
   data_col49[48] <= data_col49[47];
   data_col49[49] <= data_col49[48];

   data_col50[1] <= data[115];
   data_col50[2] <= data_col50[1];
   data_col50[3] <= data_col50[2];
   data_col50[4] <= data_col50[3];
   data_col50[5] <= data_col50[4];
   data_col50[6] <= data_col50[5];
   data_col50[7] <= data_col50[6];
   data_col50[8] <= data_col50[7];
   data_col50[9] <= data_col50[8];
   data_col50[10] <= data_col50[9];
   data_col50[11] <= data_col50[10];
   data_col50[12] <= data_col50[11];
   data_col50[13] <= data_col50[12];
   data_col50[14] <= data_col50[13];
   data_col50[15] <= data_col50[14];
   data_col50[16] <= data_col50[15];
   data_col50[17] <= data_col50[16];
   data_col50[18] <= data_col50[17];
   data_col50[19] <= data_col50[18];
   data_col50[20] <= data_col50[19];
   data_col50[21] <= data_col50[20];
   data_col50[22] <= data_col50[21];
   data_col50[23] <= data_col50[22];
   data_col50[24] <= data_col50[23];
   data_col50[25] <= data_col50[24];
   data_col50[26] <= data_col50[25];
   data_col50[27] <= data_col50[26];
   data_col50[28] <= data_col50[27];
   data_col50[29] <= data_col50[28];
   data_col50[30] <= data_col50[29];
   data_col50[31] <= data_col50[30];
   data_col50[32] <= data_col50[31];
   data_col50[33] <= data_col50[32];
   data_col50[34] <= data_col50[33];
   data_col50[35] <= data_col50[34];
   data_col50[36] <= data_col50[35];
   data_col50[37] <= data_col50[36];
   data_col50[38] <= data_col50[37];
   data_col50[39] <= data_col50[38];
   data_col50[40] <= data_col50[39];
   data_col50[41] <= data_col50[40];
   data_col50[42] <= data_col50[41];
   data_col50[43] <= data_col50[42];
   data_col50[44] <= data_col50[43];
   data_col50[45] <= data_col50[44];
   data_col50[46] <= data_col50[45];
   data_col50[47] <= data_col50[46];
   data_col50[48] <= data_col50[47];
   data_col50[49] <= data_col50[48];
   data_col50[50] <= data_col50[49];

   data_col51[1] <= data[114];
   data_col51[2] <= data_col51[1];
   data_col51[3] <= data_col51[2];
   data_col51[4] <= data_col51[3];
   data_col51[5] <= data_col51[4];
   data_col51[6] <= data_col51[5];
   data_col51[7] <= data_col51[6];
   data_col51[8] <= data_col51[7];
   data_col51[9] <= data_col51[8];
   data_col51[10] <= data_col51[9];
   data_col51[11] <= data_col51[10];
   data_col51[12] <= data_col51[11];
   data_col51[13] <= data_col51[12];
   data_col51[14] <= data_col51[13];
   data_col51[15] <= data_col51[14];
   data_col51[16] <= data_col51[15];
   data_col51[17] <= data_col51[16];
   data_col51[18] <= data_col51[17];
   data_col51[19] <= data_col51[18];
   data_col51[20] <= data_col51[19];
   data_col51[21] <= data_col51[20];
   data_col51[22] <= data_col51[21];
   data_col51[23] <= data_col51[22];
   data_col51[24] <= data_col51[23];
   data_col51[25] <= data_col51[24];
   data_col51[26] <= data_col51[25];
   data_col51[27] <= data_col51[26];
   data_col51[28] <= data_col51[27];
   data_col51[29] <= data_col51[28];
   data_col51[30] <= data_col51[29];
   data_col51[31] <= data_col51[30];
   data_col51[32] <= data_col51[31];
   data_col51[33] <= data_col51[32];
   data_col51[34] <= data_col51[33];
   data_col51[35] <= data_col51[34];
   data_col51[36] <= data_col51[35];
   data_col51[37] <= data_col51[36];
   data_col51[38] <= data_col51[37];
   data_col51[39] <= data_col51[38];
   data_col51[40] <= data_col51[39];
   data_col51[41] <= data_col51[40];
   data_col51[42] <= data_col51[41];
   data_col51[43] <= data_col51[42];
   data_col51[44] <= data_col51[43];
   data_col51[45] <= data_col51[44];
   data_col51[46] <= data_col51[45];
   data_col51[47] <= data_col51[46];
   data_col51[48] <= data_col51[47];
   data_col51[49] <= data_col51[48];
   data_col51[50] <= data_col51[49];
   data_col51[51] <= data_col51[50];

   data_col52[1] <= data[113];
   data_col52[2] <= data_col52[1];
   data_col52[3] <= data_col52[2];
   data_col52[4] <= data_col52[3];
   data_col52[5] <= data_col52[4];
   data_col52[6] <= data_col52[5];
   data_col52[7] <= data_col52[6];
   data_col52[8] <= data_col52[7];
   data_col52[9] <= data_col52[8];
   data_col52[10] <= data_col52[9];
   data_col52[11] <= data_col52[10];
   data_col52[12] <= data_col52[11];
   data_col52[13] <= data_col52[12];
   data_col52[14] <= data_col52[13];
   data_col52[15] <= data_col52[14];
   data_col52[16] <= data_col52[15];
   data_col52[17] <= data_col52[16];
   data_col52[18] <= data_col52[17];
   data_col52[19] <= data_col52[18];
   data_col52[20] <= data_col52[19];
   data_col52[21] <= data_col52[20];
   data_col52[22] <= data_col52[21];
   data_col52[23] <= data_col52[22];
   data_col52[24] <= data_col52[23];
   data_col52[25] <= data_col52[24];
   data_col52[26] <= data_col52[25];
   data_col52[27] <= data_col52[26];
   data_col52[28] <= data_col52[27];
   data_col52[29] <= data_col52[28];
   data_col52[30] <= data_col52[29];
   data_col52[31] <= data_col52[30];
   data_col52[32] <= data_col52[31];
   data_col52[33] <= data_col52[32];
   data_col52[34] <= data_col52[33];
   data_col52[35] <= data_col52[34];
   data_col52[36] <= data_col52[35];
   data_col52[37] <= data_col52[36];
   data_col52[38] <= data_col52[37];
   data_col52[39] <= data_col52[38];
   data_col52[40] <= data_col52[39];
   data_col52[41] <= data_col52[40];
   data_col52[42] <= data_col52[41];
   data_col52[43] <= data_col52[42];
   data_col52[44] <= data_col52[43];
   data_col52[45] <= data_col52[44];
   data_col52[46] <= data_col52[45];
   data_col52[47] <= data_col52[46];
   data_col52[48] <= data_col52[47];
   data_col52[49] <= data_col52[48];
   data_col52[50] <= data_col52[49];
   data_col52[51] <= data_col52[50];
   data_col52[52] <= data_col52[51];

   data_col53[1] <= data[112];
   data_col53[2] <= data_col53[1];
   data_col53[3] <= data_col53[2];
   data_col53[4] <= data_col53[3];
   data_col53[5] <= data_col53[4];
   data_col53[6] <= data_col53[5];
   data_col53[7] <= data_col53[6];
   data_col53[8] <= data_col53[7];
   data_col53[9] <= data_col53[8];
   data_col53[10] <= data_col53[9];
   data_col53[11] <= data_col53[10];
   data_col53[12] <= data_col53[11];
   data_col53[13] <= data_col53[12];
   data_col53[14] <= data_col53[13];
   data_col53[15] <= data_col53[14];
   data_col53[16] <= data_col53[15];
   data_col53[17] <= data_col53[16];
   data_col53[18] <= data_col53[17];
   data_col53[19] <= data_col53[18];
   data_col53[20] <= data_col53[19];
   data_col53[21] <= data_col53[20];
   data_col53[22] <= data_col53[21];
   data_col53[23] <= data_col53[22];
   data_col53[24] <= data_col53[23];
   data_col53[25] <= data_col53[24];
   data_col53[26] <= data_col53[25];
   data_col53[27] <= data_col53[26];
   data_col53[28] <= data_col53[27];
   data_col53[29] <= data_col53[28];
   data_col53[30] <= data_col53[29];
   data_col53[31] <= data_col53[30];
   data_col53[32] <= data_col53[31];
   data_col53[33] <= data_col53[32];
   data_col53[34] <= data_col53[33];
   data_col53[35] <= data_col53[34];
   data_col53[36] <= data_col53[35];
   data_col53[37] <= data_col53[36];
   data_col53[38] <= data_col53[37];
   data_col53[39] <= data_col53[38];
   data_col53[40] <= data_col53[39];
   data_col53[41] <= data_col53[40];
   data_col53[42] <= data_col53[41];
   data_col53[43] <= data_col53[42];
   data_col53[44] <= data_col53[43];
   data_col53[45] <= data_col53[44];
   data_col53[46] <= data_col53[45];
   data_col53[47] <= data_col53[46];
   data_col53[48] <= data_col53[47];
   data_col53[49] <= data_col53[48];
   data_col53[50] <= data_col53[49];
   data_col53[51] <= data_col53[50];
   data_col53[52] <= data_col53[51];
   data_col53[53] <= data_col53[52];

   data_col54[1] <= data[111];
   data_col54[2] <= data_col54[1];
   data_col54[3] <= data_col54[2];
   data_col54[4] <= data_col54[3];
   data_col54[5] <= data_col54[4];
   data_col54[6] <= data_col54[5];
   data_col54[7] <= data_col54[6];
   data_col54[8] <= data_col54[7];
   data_col54[9] <= data_col54[8];
   data_col54[10] <= data_col54[9];
   data_col54[11] <= data_col54[10];
   data_col54[12] <= data_col54[11];
   data_col54[13] <= data_col54[12];
   data_col54[14] <= data_col54[13];
   data_col54[15] <= data_col54[14];
   data_col54[16] <= data_col54[15];
   data_col54[17] <= data_col54[16];
   data_col54[18] <= data_col54[17];
   data_col54[19] <= data_col54[18];
   data_col54[20] <= data_col54[19];
   data_col54[21] <= data_col54[20];
   data_col54[22] <= data_col54[21];
   data_col54[23] <= data_col54[22];
   data_col54[24] <= data_col54[23];
   data_col54[25] <= data_col54[24];
   data_col54[26] <= data_col54[25];
   data_col54[27] <= data_col54[26];
   data_col54[28] <= data_col54[27];
   data_col54[29] <= data_col54[28];
   data_col54[30] <= data_col54[29];
   data_col54[31] <= data_col54[30];
   data_col54[32] <= data_col54[31];
   data_col54[33] <= data_col54[32];
   data_col54[34] <= data_col54[33];
   data_col54[35] <= data_col54[34];
   data_col54[36] <= data_col54[35];
   data_col54[37] <= data_col54[36];
   data_col54[38] <= data_col54[37];
   data_col54[39] <= data_col54[38];
   data_col54[40] <= data_col54[39];
   data_col54[41] <= data_col54[40];
   data_col54[42] <= data_col54[41];
   data_col54[43] <= data_col54[42];
   data_col54[44] <= data_col54[43];
   data_col54[45] <= data_col54[44];
   data_col54[46] <= data_col54[45];
   data_col54[47] <= data_col54[46];
   data_col54[48] <= data_col54[47];
   data_col54[49] <= data_col54[48];
   data_col54[50] <= data_col54[49];
   data_col54[51] <= data_col54[50];
   data_col54[52] <= data_col54[51];
   data_col54[53] <= data_col54[52];
   data_col54[54] <= data_col54[53];

   data_col55[1] <= data[110];
   data_col55[2] <= data_col55[1];
   data_col55[3] <= data_col55[2];
   data_col55[4] <= data_col55[3];
   data_col55[5] <= data_col55[4];
   data_col55[6] <= data_col55[5];
   data_col55[7] <= data_col55[6];
   data_col55[8] <= data_col55[7];
   data_col55[9] <= data_col55[8];
   data_col55[10] <= data_col55[9];
   data_col55[11] <= data_col55[10];
   data_col55[12] <= data_col55[11];
   data_col55[13] <= data_col55[12];
   data_col55[14] <= data_col55[13];
   data_col55[15] <= data_col55[14];
   data_col55[16] <= data_col55[15];
   data_col55[17] <= data_col55[16];
   data_col55[18] <= data_col55[17];
   data_col55[19] <= data_col55[18];
   data_col55[20] <= data_col55[19];
   data_col55[21] <= data_col55[20];
   data_col55[22] <= data_col55[21];
   data_col55[23] <= data_col55[22];
   data_col55[24] <= data_col55[23];
   data_col55[25] <= data_col55[24];
   data_col55[26] <= data_col55[25];
   data_col55[27] <= data_col55[26];
   data_col55[28] <= data_col55[27];
   data_col55[29] <= data_col55[28];
   data_col55[30] <= data_col55[29];
   data_col55[31] <= data_col55[30];
   data_col55[32] <= data_col55[31];
   data_col55[33] <= data_col55[32];
   data_col55[34] <= data_col55[33];
   data_col55[35] <= data_col55[34];
   data_col55[36] <= data_col55[35];
   data_col55[37] <= data_col55[36];
   data_col55[38] <= data_col55[37];
   data_col55[39] <= data_col55[38];
   data_col55[40] <= data_col55[39];
   data_col55[41] <= data_col55[40];
   data_col55[42] <= data_col55[41];
   data_col55[43] <= data_col55[42];
   data_col55[44] <= data_col55[43];
   data_col55[45] <= data_col55[44];
   data_col55[46] <= data_col55[45];
   data_col55[47] <= data_col55[46];
   data_col55[48] <= data_col55[47];
   data_col55[49] <= data_col55[48];
   data_col55[50] <= data_col55[49];
   data_col55[51] <= data_col55[50];
   data_col55[52] <= data_col55[51];
   data_col55[53] <= data_col55[52];
   data_col55[54] <= data_col55[53];
   data_col55[55] <= data_col55[54];

   data_col56[1] <= data[109];
   data_col56[2] <= data_col56[1];
   data_col56[3] <= data_col56[2];
   data_col56[4] <= data_col56[3];
   data_col56[5] <= data_col56[4];
   data_col56[6] <= data_col56[5];
   data_col56[7] <= data_col56[6];
   data_col56[8] <= data_col56[7];
   data_col56[9] <= data_col56[8];
   data_col56[10] <= data_col56[9];
   data_col56[11] <= data_col56[10];
   data_col56[12] <= data_col56[11];
   data_col56[13] <= data_col56[12];
   data_col56[14] <= data_col56[13];
   data_col56[15] <= data_col56[14];
   data_col56[16] <= data_col56[15];
   data_col56[17] <= data_col56[16];
   data_col56[18] <= data_col56[17];
   data_col56[19] <= data_col56[18];
   data_col56[20] <= data_col56[19];
   data_col56[21] <= data_col56[20];
   data_col56[22] <= data_col56[21];
   data_col56[23] <= data_col56[22];
   data_col56[24] <= data_col56[23];
   data_col56[25] <= data_col56[24];
   data_col56[26] <= data_col56[25];
   data_col56[27] <= data_col56[26];
   data_col56[28] <= data_col56[27];
   data_col56[29] <= data_col56[28];
   data_col56[30] <= data_col56[29];
   data_col56[31] <= data_col56[30];
   data_col56[32] <= data_col56[31];
   data_col56[33] <= data_col56[32];
   data_col56[34] <= data_col56[33];
   data_col56[35] <= data_col56[34];
   data_col56[36] <= data_col56[35];
   data_col56[37] <= data_col56[36];
   data_col56[38] <= data_col56[37];
   data_col56[39] <= data_col56[38];
   data_col56[40] <= data_col56[39];
   data_col56[41] <= data_col56[40];
   data_col56[42] <= data_col56[41];
   data_col56[43] <= data_col56[42];
   data_col56[44] <= data_col56[43];
   data_col56[45] <= data_col56[44];
   data_col56[46] <= data_col56[45];
   data_col56[47] <= data_col56[46];
   data_col56[48] <= data_col56[47];
   data_col56[49] <= data_col56[48];
   data_col56[50] <= data_col56[49];
   data_col56[51] <= data_col56[50];
   data_col56[52] <= data_col56[51];
   data_col56[53] <= data_col56[52];
   data_col56[54] <= data_col56[53];
   data_col56[55] <= data_col56[54];
   data_col56[56] <= data_col56[55];

   data_col57[1] <= data[108];
   data_col57[2] <= data_col57[1];
   data_col57[3] <= data_col57[2];
   data_col57[4] <= data_col57[3];
   data_col57[5] <= data_col57[4];
   data_col57[6] <= data_col57[5];
   data_col57[7] <= data_col57[6];
   data_col57[8] <= data_col57[7];
   data_col57[9] <= data_col57[8];
   data_col57[10] <= data_col57[9];
   data_col57[11] <= data_col57[10];
   data_col57[12] <= data_col57[11];
   data_col57[13] <= data_col57[12];
   data_col57[14] <= data_col57[13];
   data_col57[15] <= data_col57[14];
   data_col57[16] <= data_col57[15];
   data_col57[17] <= data_col57[16];
   data_col57[18] <= data_col57[17];
   data_col57[19] <= data_col57[18];
   data_col57[20] <= data_col57[19];
   data_col57[21] <= data_col57[20];
   data_col57[22] <= data_col57[21];
   data_col57[23] <= data_col57[22];
   data_col57[24] <= data_col57[23];
   data_col57[25] <= data_col57[24];
   data_col57[26] <= data_col57[25];
   data_col57[27] <= data_col57[26];
   data_col57[28] <= data_col57[27];
   data_col57[29] <= data_col57[28];
   data_col57[30] <= data_col57[29];
   data_col57[31] <= data_col57[30];
   data_col57[32] <= data_col57[31];
   data_col57[33] <= data_col57[32];
   data_col57[34] <= data_col57[33];
   data_col57[35] <= data_col57[34];
   data_col57[36] <= data_col57[35];
   data_col57[37] <= data_col57[36];
   data_col57[38] <= data_col57[37];
   data_col57[39] <= data_col57[38];
   data_col57[40] <= data_col57[39];
   data_col57[41] <= data_col57[40];
   data_col57[42] <= data_col57[41];
   data_col57[43] <= data_col57[42];
   data_col57[44] <= data_col57[43];
   data_col57[45] <= data_col57[44];
   data_col57[46] <= data_col57[45];
   data_col57[47] <= data_col57[46];
   data_col57[48] <= data_col57[47];
   data_col57[49] <= data_col57[48];
   data_col57[50] <= data_col57[49];
   data_col57[51] <= data_col57[50];
   data_col57[52] <= data_col57[51];
   data_col57[53] <= data_col57[52];
   data_col57[54] <= data_col57[53];
   data_col57[55] <= data_col57[54];
   data_col57[56] <= data_col57[55];
   data_col57[57] <= data_col57[56];

   data_col58[1] <= data[107];
   data_col58[2] <= data_col58[1];
   data_col58[3] <= data_col58[2];
   data_col58[4] <= data_col58[3];
   data_col58[5] <= data_col58[4];
   data_col58[6] <= data_col58[5];
   data_col58[7] <= data_col58[6];
   data_col58[8] <= data_col58[7];
   data_col58[9] <= data_col58[8];
   data_col58[10] <= data_col58[9];
   data_col58[11] <= data_col58[10];
   data_col58[12] <= data_col58[11];
   data_col58[13] <= data_col58[12];
   data_col58[14] <= data_col58[13];
   data_col58[15] <= data_col58[14];
   data_col58[16] <= data_col58[15];
   data_col58[17] <= data_col58[16];
   data_col58[18] <= data_col58[17];
   data_col58[19] <= data_col58[18];
   data_col58[20] <= data_col58[19];
   data_col58[21] <= data_col58[20];
   data_col58[22] <= data_col58[21];
   data_col58[23] <= data_col58[22];
   data_col58[24] <= data_col58[23];
   data_col58[25] <= data_col58[24];
   data_col58[26] <= data_col58[25];
   data_col58[27] <= data_col58[26];
   data_col58[28] <= data_col58[27];
   data_col58[29] <= data_col58[28];
   data_col58[30] <= data_col58[29];
   data_col58[31] <= data_col58[30];
   data_col58[32] <= data_col58[31];
   data_col58[33] <= data_col58[32];
   data_col58[34] <= data_col58[33];
   data_col58[35] <= data_col58[34];
   data_col58[36] <= data_col58[35];
   data_col58[37] <= data_col58[36];
   data_col58[38] <= data_col58[37];
   data_col58[39] <= data_col58[38];
   data_col58[40] <= data_col58[39];
   data_col58[41] <= data_col58[40];
   data_col58[42] <= data_col58[41];
   data_col58[43] <= data_col58[42];
   data_col58[44] <= data_col58[43];
   data_col58[45] <= data_col58[44];
   data_col58[46] <= data_col58[45];
   data_col58[47] <= data_col58[46];
   data_col58[48] <= data_col58[47];
   data_col58[49] <= data_col58[48];
   data_col58[50] <= data_col58[49];
   data_col58[51] <= data_col58[50];
   data_col58[52] <= data_col58[51];
   data_col58[53] <= data_col58[52];
   data_col58[54] <= data_col58[53];
   data_col58[55] <= data_col58[54];
   data_col58[56] <= data_col58[55];
   data_col58[57] <= data_col58[56];
   data_col58[58] <= data_col58[57];

   data_col59[1] <= data[106];
   data_col59[2] <= data_col59[1];
   data_col59[3] <= data_col59[2];
   data_col59[4] <= data_col59[3];
   data_col59[5] <= data_col59[4];
   data_col59[6] <= data_col59[5];
   data_col59[7] <= data_col59[6];
   data_col59[8] <= data_col59[7];
   data_col59[9] <= data_col59[8];
   data_col59[10] <= data_col59[9];
   data_col59[11] <= data_col59[10];
   data_col59[12] <= data_col59[11];
   data_col59[13] <= data_col59[12];
   data_col59[14] <= data_col59[13];
   data_col59[15] <= data_col59[14];
   data_col59[16] <= data_col59[15];
   data_col59[17] <= data_col59[16];
   data_col59[18] <= data_col59[17];
   data_col59[19] <= data_col59[18];
   data_col59[20] <= data_col59[19];
   data_col59[21] <= data_col59[20];
   data_col59[22] <= data_col59[21];
   data_col59[23] <= data_col59[22];
   data_col59[24] <= data_col59[23];
   data_col59[25] <= data_col59[24];
   data_col59[26] <= data_col59[25];
   data_col59[27] <= data_col59[26];
   data_col59[28] <= data_col59[27];
   data_col59[29] <= data_col59[28];
   data_col59[30] <= data_col59[29];
   data_col59[31] <= data_col59[30];
   data_col59[32] <= data_col59[31];
   data_col59[33] <= data_col59[32];
   data_col59[34] <= data_col59[33];
   data_col59[35] <= data_col59[34];
   data_col59[36] <= data_col59[35];
   data_col59[37] <= data_col59[36];
   data_col59[38] <= data_col59[37];
   data_col59[39] <= data_col59[38];
   data_col59[40] <= data_col59[39];
   data_col59[41] <= data_col59[40];
   data_col59[42] <= data_col59[41];
   data_col59[43] <= data_col59[42];
   data_col59[44] <= data_col59[43];
   data_col59[45] <= data_col59[44];
   data_col59[46] <= data_col59[45];
   data_col59[47] <= data_col59[46];
   data_col59[48] <= data_col59[47];
   data_col59[49] <= data_col59[48];
   data_col59[50] <= data_col59[49];
   data_col59[51] <= data_col59[50];
   data_col59[52] <= data_col59[51];
   data_col59[53] <= data_col59[52];
   data_col59[54] <= data_col59[53];
   data_col59[55] <= data_col59[54];
   data_col59[56] <= data_col59[55];
   data_col59[57] <= data_col59[56];
   data_col59[58] <= data_col59[57];
   data_col59[59] <= data_col59[58];

   data_col60[1] <= data[105];
   data_col60[2] <= data_col60[1];
   data_col60[3] <= data_col60[2];
   data_col60[4] <= data_col60[3];
   data_col60[5] <= data_col60[4];
   data_col60[6] <= data_col60[5];
   data_col60[7] <= data_col60[6];
   data_col60[8] <= data_col60[7];
   data_col60[9] <= data_col60[8];
   data_col60[10] <= data_col60[9];
   data_col60[11] <= data_col60[10];
   data_col60[12] <= data_col60[11];
   data_col60[13] <= data_col60[12];
   data_col60[14] <= data_col60[13];
   data_col60[15] <= data_col60[14];
   data_col60[16] <= data_col60[15];
   data_col60[17] <= data_col60[16];
   data_col60[18] <= data_col60[17];
   data_col60[19] <= data_col60[18];
   data_col60[20] <= data_col60[19];
   data_col60[21] <= data_col60[20];
   data_col60[22] <= data_col60[21];
   data_col60[23] <= data_col60[22];
   data_col60[24] <= data_col60[23];
   data_col60[25] <= data_col60[24];
   data_col60[26] <= data_col60[25];
   data_col60[27] <= data_col60[26];
   data_col60[28] <= data_col60[27];
   data_col60[29] <= data_col60[28];
   data_col60[30] <= data_col60[29];
   data_col60[31] <= data_col60[30];
   data_col60[32] <= data_col60[31];
   data_col60[33] <= data_col60[32];
   data_col60[34] <= data_col60[33];
   data_col60[35] <= data_col60[34];
   data_col60[36] <= data_col60[35];
   data_col60[37] <= data_col60[36];
   data_col60[38] <= data_col60[37];
   data_col60[39] <= data_col60[38];
   data_col60[40] <= data_col60[39];
   data_col60[41] <= data_col60[40];
   data_col60[42] <= data_col60[41];
   data_col60[43] <= data_col60[42];
   data_col60[44] <= data_col60[43];
   data_col60[45] <= data_col60[44];
   data_col60[46] <= data_col60[45];
   data_col60[47] <= data_col60[46];
   data_col60[48] <= data_col60[47];
   data_col60[49] <= data_col60[48];
   data_col60[50] <= data_col60[49];
   data_col60[51] <= data_col60[50];
   data_col60[52] <= data_col60[51];
   data_col60[53] <= data_col60[52];
   data_col60[54] <= data_col60[53];
   data_col60[55] <= data_col60[54];
   data_col60[56] <= data_col60[55];
   data_col60[57] <= data_col60[56];
   data_col60[58] <= data_col60[57];
   data_col60[59] <= data_col60[58];
   data_col60[60] <= data_col60[59];

   data_col61[1] <= data[104];
   data_col61[2] <= data_col61[1];
   data_col61[3] <= data_col61[2];
   data_col61[4] <= data_col61[3];
   data_col61[5] <= data_col61[4];
   data_col61[6] <= data_col61[5];
   data_col61[7] <= data_col61[6];
   data_col61[8] <= data_col61[7];
   data_col61[9] <= data_col61[8];
   data_col61[10] <= data_col61[9];
   data_col61[11] <= data_col61[10];
   data_col61[12] <= data_col61[11];
   data_col61[13] <= data_col61[12];
   data_col61[14] <= data_col61[13];
   data_col61[15] <= data_col61[14];
   data_col61[16] <= data_col61[15];
   data_col61[17] <= data_col61[16];
   data_col61[18] <= data_col61[17];
   data_col61[19] <= data_col61[18];
   data_col61[20] <= data_col61[19];
   data_col61[21] <= data_col61[20];
   data_col61[22] <= data_col61[21];
   data_col61[23] <= data_col61[22];
   data_col61[24] <= data_col61[23];
   data_col61[25] <= data_col61[24];
   data_col61[26] <= data_col61[25];
   data_col61[27] <= data_col61[26];
   data_col61[28] <= data_col61[27];
   data_col61[29] <= data_col61[28];
   data_col61[30] <= data_col61[29];
   data_col61[31] <= data_col61[30];
   data_col61[32] <= data_col61[31];
   data_col61[33] <= data_col61[32];
   data_col61[34] <= data_col61[33];
   data_col61[35] <= data_col61[34];
   data_col61[36] <= data_col61[35];
   data_col61[37] <= data_col61[36];
   data_col61[38] <= data_col61[37];
   data_col61[39] <= data_col61[38];
   data_col61[40] <= data_col61[39];
   data_col61[41] <= data_col61[40];
   data_col61[42] <= data_col61[41];
   data_col61[43] <= data_col61[42];
   data_col61[44] <= data_col61[43];
   data_col61[45] <= data_col61[44];
   data_col61[46] <= data_col61[45];
   data_col61[47] <= data_col61[46];
   data_col61[48] <= data_col61[47];
   data_col61[49] <= data_col61[48];
   data_col61[50] <= data_col61[49];
   data_col61[51] <= data_col61[50];
   data_col61[52] <= data_col61[51];
   data_col61[53] <= data_col61[52];
   data_col61[54] <= data_col61[53];
   data_col61[55] <= data_col61[54];
   data_col61[56] <= data_col61[55];
   data_col61[57] <= data_col61[56];
   data_col61[58] <= data_col61[57];
   data_col61[59] <= data_col61[58];
   data_col61[60] <= data_col61[59];
   data_col61[61] <= data_col61[60];

   data_col62[1] <= data[103];
   data_col62[2] <= data_col62[1];
   data_col62[3] <= data_col62[2];
   data_col62[4] <= data_col62[3];
   data_col62[5] <= data_col62[4];
   data_col62[6] <= data_col62[5];
   data_col62[7] <= data_col62[6];
   data_col62[8] <= data_col62[7];
   data_col62[9] <= data_col62[8];
   data_col62[10] <= data_col62[9];
   data_col62[11] <= data_col62[10];
   data_col62[12] <= data_col62[11];
   data_col62[13] <= data_col62[12];
   data_col62[14] <= data_col62[13];
   data_col62[15] <= data_col62[14];
   data_col62[16] <= data_col62[15];
   data_col62[17] <= data_col62[16];
   data_col62[18] <= data_col62[17];
   data_col62[19] <= data_col62[18];
   data_col62[20] <= data_col62[19];
   data_col62[21] <= data_col62[20];
   data_col62[22] <= data_col62[21];
   data_col62[23] <= data_col62[22];
   data_col62[24] <= data_col62[23];
   data_col62[25] <= data_col62[24];
   data_col62[26] <= data_col62[25];
   data_col62[27] <= data_col62[26];
   data_col62[28] <= data_col62[27];
   data_col62[29] <= data_col62[28];
   data_col62[30] <= data_col62[29];
   data_col62[31] <= data_col62[30];
   data_col62[32] <= data_col62[31];
   data_col62[33] <= data_col62[32];
   data_col62[34] <= data_col62[33];
   data_col62[35] <= data_col62[34];
   data_col62[36] <= data_col62[35];
   data_col62[37] <= data_col62[36];
   data_col62[38] <= data_col62[37];
   data_col62[39] <= data_col62[38];
   data_col62[40] <= data_col62[39];
   data_col62[41] <= data_col62[40];
   data_col62[42] <= data_col62[41];
   data_col62[43] <= data_col62[42];
   data_col62[44] <= data_col62[43];
   data_col62[45] <= data_col62[44];
   data_col62[46] <= data_col62[45];
   data_col62[47] <= data_col62[46];
   data_col62[48] <= data_col62[47];
   data_col62[49] <= data_col62[48];
   data_col62[50] <= data_col62[49];
   data_col62[51] <= data_col62[50];
   data_col62[52] <= data_col62[51];
   data_col62[53] <= data_col62[52];
   data_col62[54] <= data_col62[53];
   data_col62[55] <= data_col62[54];
   data_col62[56] <= data_col62[55];
   data_col62[57] <= data_col62[56];
   data_col62[58] <= data_col62[57];
   data_col62[59] <= data_col62[58];
   data_col62[60] <= data_col62[59];
   data_col62[61] <= data_col62[60];
   data_col62[62] <= data_col62[61];

   data_col63[1] <= data[102];
   data_col63[2] <= data_col63[1];
   data_col63[3] <= data_col63[2];
   data_col63[4] <= data_col63[3];
   data_col63[5] <= data_col63[4];
   data_col63[6] <= data_col63[5];
   data_col63[7] <= data_col63[6];
   data_col63[8] <= data_col63[7];
   data_col63[9] <= data_col63[8];
   data_col63[10] <= data_col63[9];
   data_col63[11] <= data_col63[10];
   data_col63[12] <= data_col63[11];
   data_col63[13] <= data_col63[12];
   data_col63[14] <= data_col63[13];
   data_col63[15] <= data_col63[14];
   data_col63[16] <= data_col63[15];
   data_col63[17] <= data_col63[16];
   data_col63[18] <= data_col63[17];
   data_col63[19] <= data_col63[18];
   data_col63[20] <= data_col63[19];
   data_col63[21] <= data_col63[20];
   data_col63[22] <= data_col63[21];
   data_col63[23] <= data_col63[22];
   data_col63[24] <= data_col63[23];
   data_col63[25] <= data_col63[24];
   data_col63[26] <= data_col63[25];
   data_col63[27] <= data_col63[26];
   data_col63[28] <= data_col63[27];
   data_col63[29] <= data_col63[28];
   data_col63[30] <= data_col63[29];
   data_col63[31] <= data_col63[30];
   data_col63[32] <= data_col63[31];
   data_col63[33] <= data_col63[32];
   data_col63[34] <= data_col63[33];
   data_col63[35] <= data_col63[34];
   data_col63[36] <= data_col63[35];
   data_col63[37] <= data_col63[36];
   data_col63[38] <= data_col63[37];
   data_col63[39] <= data_col63[38];
   data_col63[40] <= data_col63[39];
   data_col63[41] <= data_col63[40];
   data_col63[42] <= data_col63[41];
   data_col63[43] <= data_col63[42];
   data_col63[44] <= data_col63[43];
   data_col63[45] <= data_col63[44];
   data_col63[46] <= data_col63[45];
   data_col63[47] <= data_col63[46];
   data_col63[48] <= data_col63[47];
   data_col63[49] <= data_col63[48];
   data_col63[50] <= data_col63[49];
   data_col63[51] <= data_col63[50];
   data_col63[52] <= data_col63[51];
   data_col63[53] <= data_col63[52];
   data_col63[54] <= data_col63[53];
   data_col63[55] <= data_col63[54];
   data_col63[56] <= data_col63[55];
   data_col63[57] <= data_col63[56];
   data_col63[58] <= data_col63[57];
   data_col63[59] <= data_col63[58];
   data_col63[60] <= data_col63[59];
   data_col63[61] <= data_col63[60];
   data_col63[62] <= data_col63[61];
   data_col63[63] <= data_col63[62];

   data_col64[1] <= data[101];
   data_col64[2] <= data_col64[1];
   data_col64[3] <= data_col64[2];
   data_col64[4] <= data_col64[3];
   data_col64[5] <= data_col64[4];
   data_col64[6] <= data_col64[5];
   data_col64[7] <= data_col64[6];
   data_col64[8] <= data_col64[7];
   data_col64[9] <= data_col64[8];
   data_col64[10] <= data_col64[9];
   data_col64[11] <= data_col64[10];
   data_col64[12] <= data_col64[11];
   data_col64[13] <= data_col64[12];
   data_col64[14] <= data_col64[13];
   data_col64[15] <= data_col64[14];
   data_col64[16] <= data_col64[15];
   data_col64[17] <= data_col64[16];
   data_col64[18] <= data_col64[17];
   data_col64[19] <= data_col64[18];
   data_col64[20] <= data_col64[19];
   data_col64[21] <= data_col64[20];
   data_col64[22] <= data_col64[21];
   data_col64[23] <= data_col64[22];
   data_col64[24] <= data_col64[23];
   data_col64[25] <= data_col64[24];
   data_col64[26] <= data_col64[25];
   data_col64[27] <= data_col64[26];
   data_col64[28] <= data_col64[27];
   data_col64[29] <= data_col64[28];
   data_col64[30] <= data_col64[29];
   data_col64[31] <= data_col64[30];
   data_col64[32] <= data_col64[31];
   data_col64[33] <= data_col64[32];
   data_col64[34] <= data_col64[33];
   data_col64[35] <= data_col64[34];
   data_col64[36] <= data_col64[35];
   data_col64[37] <= data_col64[36];
   data_col64[38] <= data_col64[37];
   data_col64[39] <= data_col64[38];
   data_col64[40] <= data_col64[39];
   data_col64[41] <= data_col64[40];
   data_col64[42] <= data_col64[41];
   data_col64[43] <= data_col64[42];
   data_col64[44] <= data_col64[43];
   data_col64[45] <= data_col64[44];
   data_col64[46] <= data_col64[45];
   data_col64[47] <= data_col64[46];
   data_col64[48] <= data_col64[47];
   data_col64[49] <= data_col64[48];
   data_col64[50] <= data_col64[49];
   data_col64[51] <= data_col64[50];
   data_col64[52] <= data_col64[51];
   data_col64[53] <= data_col64[52];
   data_col64[54] <= data_col64[53];
   data_col64[55] <= data_col64[54];
   data_col64[56] <= data_col64[55];
   data_col64[57] <= data_col64[56];
   data_col64[58] <= data_col64[57];
   data_col64[59] <= data_col64[58];
   data_col64[60] <= data_col64[59];
   data_col64[61] <= data_col64[60];
   data_col64[62] <= data_col64[61];
   data_col64[63] <= data_col64[62];
   data_col64[64] <= data_col64[63];

   data_col65[1] <= data[100];
   data_col65[2] <= data_col65[1];
   data_col65[3] <= data_col65[2];
   data_col65[4] <= data_col65[3];
   data_col65[5] <= data_col65[4];
   data_col65[6] <= data_col65[5];
   data_col65[7] <= data_col65[6];
   data_col65[8] <= data_col65[7];
   data_col65[9] <= data_col65[8];
   data_col65[10] <= data_col65[9];
   data_col65[11] <= data_col65[10];
   data_col65[12] <= data_col65[11];
   data_col65[13] <= data_col65[12];
   data_col65[14] <= data_col65[13];
   data_col65[15] <= data_col65[14];
   data_col65[16] <= data_col65[15];
   data_col65[17] <= data_col65[16];
   data_col65[18] <= data_col65[17];
   data_col65[19] <= data_col65[18];
   data_col65[20] <= data_col65[19];
   data_col65[21] <= data_col65[20];
   data_col65[22] <= data_col65[21];
   data_col65[23] <= data_col65[22];
   data_col65[24] <= data_col65[23];
   data_col65[25] <= data_col65[24];
   data_col65[26] <= data_col65[25];
   data_col65[27] <= data_col65[26];
   data_col65[28] <= data_col65[27];
   data_col65[29] <= data_col65[28];
   data_col65[30] <= data_col65[29];
   data_col65[31] <= data_col65[30];
   data_col65[32] <= data_col65[31];
   data_col65[33] <= data_col65[32];
   data_col65[34] <= data_col65[33];
   data_col65[35] <= data_col65[34];
   data_col65[36] <= data_col65[35];
   data_col65[37] <= data_col65[36];
   data_col65[38] <= data_col65[37];
   data_col65[39] <= data_col65[38];
   data_col65[40] <= data_col65[39];
   data_col65[41] <= data_col65[40];
   data_col65[42] <= data_col65[41];
   data_col65[43] <= data_col65[42];
   data_col65[44] <= data_col65[43];
   data_col65[45] <= data_col65[44];
   data_col65[46] <= data_col65[45];
   data_col65[47] <= data_col65[46];
   data_col65[48] <= data_col65[47];
   data_col65[49] <= data_col65[48];
   data_col65[50] <= data_col65[49];
   data_col65[51] <= data_col65[50];
   data_col65[52] <= data_col65[51];
   data_col65[53] <= data_col65[52];
   data_col65[54] <= data_col65[53];
   data_col65[55] <= data_col65[54];
   data_col65[56] <= data_col65[55];
   data_col65[57] <= data_col65[56];
   data_col65[58] <= data_col65[57];
   data_col65[59] <= data_col65[58];
   data_col65[60] <= data_col65[59];
   data_col65[61] <= data_col65[60];
   data_col65[62] <= data_col65[61];
   data_col65[63] <= data_col65[62];
   data_col65[64] <= data_col65[63];
   data_col65[65] <= data_col65[64];

   data_col66[1] <= data[99];
   data_col66[2] <= data_col66[1];
   data_col66[3] <= data_col66[2];
   data_col66[4] <= data_col66[3];
   data_col66[5] <= data_col66[4];
   data_col66[6] <= data_col66[5];
   data_col66[7] <= data_col66[6];
   data_col66[8] <= data_col66[7];
   data_col66[9] <= data_col66[8];
   data_col66[10] <= data_col66[9];
   data_col66[11] <= data_col66[10];
   data_col66[12] <= data_col66[11];
   data_col66[13] <= data_col66[12];
   data_col66[14] <= data_col66[13];
   data_col66[15] <= data_col66[14];
   data_col66[16] <= data_col66[15];
   data_col66[17] <= data_col66[16];
   data_col66[18] <= data_col66[17];
   data_col66[19] <= data_col66[18];
   data_col66[20] <= data_col66[19];
   data_col66[21] <= data_col66[20];
   data_col66[22] <= data_col66[21];
   data_col66[23] <= data_col66[22];
   data_col66[24] <= data_col66[23];
   data_col66[25] <= data_col66[24];
   data_col66[26] <= data_col66[25];
   data_col66[27] <= data_col66[26];
   data_col66[28] <= data_col66[27];
   data_col66[29] <= data_col66[28];
   data_col66[30] <= data_col66[29];
   data_col66[31] <= data_col66[30];
   data_col66[32] <= data_col66[31];
   data_col66[33] <= data_col66[32];
   data_col66[34] <= data_col66[33];
   data_col66[35] <= data_col66[34];
   data_col66[36] <= data_col66[35];
   data_col66[37] <= data_col66[36];
   data_col66[38] <= data_col66[37];
   data_col66[39] <= data_col66[38];
   data_col66[40] <= data_col66[39];
   data_col66[41] <= data_col66[40];
   data_col66[42] <= data_col66[41];
   data_col66[43] <= data_col66[42];
   data_col66[44] <= data_col66[43];
   data_col66[45] <= data_col66[44];
   data_col66[46] <= data_col66[45];
   data_col66[47] <= data_col66[46];
   data_col66[48] <= data_col66[47];
   data_col66[49] <= data_col66[48];
   data_col66[50] <= data_col66[49];
   data_col66[51] <= data_col66[50];
   data_col66[52] <= data_col66[51];
   data_col66[53] <= data_col66[52];
   data_col66[54] <= data_col66[53];
   data_col66[55] <= data_col66[54];
   data_col66[56] <= data_col66[55];
   data_col66[57] <= data_col66[56];
   data_col66[58] <= data_col66[57];
   data_col66[59] <= data_col66[58];
   data_col66[60] <= data_col66[59];
   data_col66[61] <= data_col66[60];
   data_col66[62] <= data_col66[61];
   data_col66[63] <= data_col66[62];
   data_col66[64] <= data_col66[63];
   data_col66[65] <= data_col66[64];
   data_col66[66] <= data_col66[65];

   data_col67[1] <= data[98];
   data_col67[2] <= data_col67[1];
   data_col67[3] <= data_col67[2];
   data_col67[4] <= data_col67[3];
   data_col67[5] <= data_col67[4];
   data_col67[6] <= data_col67[5];
   data_col67[7] <= data_col67[6];
   data_col67[8] <= data_col67[7];
   data_col67[9] <= data_col67[8];
   data_col67[10] <= data_col67[9];
   data_col67[11] <= data_col67[10];
   data_col67[12] <= data_col67[11];
   data_col67[13] <= data_col67[12];
   data_col67[14] <= data_col67[13];
   data_col67[15] <= data_col67[14];
   data_col67[16] <= data_col67[15];
   data_col67[17] <= data_col67[16];
   data_col67[18] <= data_col67[17];
   data_col67[19] <= data_col67[18];
   data_col67[20] <= data_col67[19];
   data_col67[21] <= data_col67[20];
   data_col67[22] <= data_col67[21];
   data_col67[23] <= data_col67[22];
   data_col67[24] <= data_col67[23];
   data_col67[25] <= data_col67[24];
   data_col67[26] <= data_col67[25];
   data_col67[27] <= data_col67[26];
   data_col67[28] <= data_col67[27];
   data_col67[29] <= data_col67[28];
   data_col67[30] <= data_col67[29];
   data_col67[31] <= data_col67[30];
   data_col67[32] <= data_col67[31];
   data_col67[33] <= data_col67[32];
   data_col67[34] <= data_col67[33];
   data_col67[35] <= data_col67[34];
   data_col67[36] <= data_col67[35];
   data_col67[37] <= data_col67[36];
   data_col67[38] <= data_col67[37];
   data_col67[39] <= data_col67[38];
   data_col67[40] <= data_col67[39];
   data_col67[41] <= data_col67[40];
   data_col67[42] <= data_col67[41];
   data_col67[43] <= data_col67[42];
   data_col67[44] <= data_col67[43];
   data_col67[45] <= data_col67[44];
   data_col67[46] <= data_col67[45];
   data_col67[47] <= data_col67[46];
   data_col67[48] <= data_col67[47];
   data_col67[49] <= data_col67[48];
   data_col67[50] <= data_col67[49];
   data_col67[51] <= data_col67[50];
   data_col67[52] <= data_col67[51];
   data_col67[53] <= data_col67[52];
   data_col67[54] <= data_col67[53];
   data_col67[55] <= data_col67[54];
   data_col67[56] <= data_col67[55];
   data_col67[57] <= data_col67[56];
   data_col67[58] <= data_col67[57];
   data_col67[59] <= data_col67[58];
   data_col67[60] <= data_col67[59];
   data_col67[61] <= data_col67[60];
   data_col67[62] <= data_col67[61];
   data_col67[63] <= data_col67[62];
   data_col67[64] <= data_col67[63];
   data_col67[65] <= data_col67[64];
   data_col67[66] <= data_col67[65];
   data_col67[67] <= data_col67[66];

   data_col68[1] <= data[97];
   data_col68[2] <= data_col68[1];
   data_col68[3] <= data_col68[2];
   data_col68[4] <= data_col68[3];
   data_col68[5] <= data_col68[4];
   data_col68[6] <= data_col68[5];
   data_col68[7] <= data_col68[6];
   data_col68[8] <= data_col68[7];
   data_col68[9] <= data_col68[8];
   data_col68[10] <= data_col68[9];
   data_col68[11] <= data_col68[10];
   data_col68[12] <= data_col68[11];
   data_col68[13] <= data_col68[12];
   data_col68[14] <= data_col68[13];
   data_col68[15] <= data_col68[14];
   data_col68[16] <= data_col68[15];
   data_col68[17] <= data_col68[16];
   data_col68[18] <= data_col68[17];
   data_col68[19] <= data_col68[18];
   data_col68[20] <= data_col68[19];
   data_col68[21] <= data_col68[20];
   data_col68[22] <= data_col68[21];
   data_col68[23] <= data_col68[22];
   data_col68[24] <= data_col68[23];
   data_col68[25] <= data_col68[24];
   data_col68[26] <= data_col68[25];
   data_col68[27] <= data_col68[26];
   data_col68[28] <= data_col68[27];
   data_col68[29] <= data_col68[28];
   data_col68[30] <= data_col68[29];
   data_col68[31] <= data_col68[30];
   data_col68[32] <= data_col68[31];
   data_col68[33] <= data_col68[32];
   data_col68[34] <= data_col68[33];
   data_col68[35] <= data_col68[34];
   data_col68[36] <= data_col68[35];
   data_col68[37] <= data_col68[36];
   data_col68[38] <= data_col68[37];
   data_col68[39] <= data_col68[38];
   data_col68[40] <= data_col68[39];
   data_col68[41] <= data_col68[40];
   data_col68[42] <= data_col68[41];
   data_col68[43] <= data_col68[42];
   data_col68[44] <= data_col68[43];
   data_col68[45] <= data_col68[44];
   data_col68[46] <= data_col68[45];
   data_col68[47] <= data_col68[46];
   data_col68[48] <= data_col68[47];
   data_col68[49] <= data_col68[48];
   data_col68[50] <= data_col68[49];
   data_col68[51] <= data_col68[50];
   data_col68[52] <= data_col68[51];
   data_col68[53] <= data_col68[52];
   data_col68[54] <= data_col68[53];
   data_col68[55] <= data_col68[54];
   data_col68[56] <= data_col68[55];
   data_col68[57] <= data_col68[56];
   data_col68[58] <= data_col68[57];
   data_col68[59] <= data_col68[58];
   data_col68[60] <= data_col68[59];
   data_col68[61] <= data_col68[60];
   data_col68[62] <= data_col68[61];
   data_col68[63] <= data_col68[62];
   data_col68[64] <= data_col68[63];
   data_col68[65] <= data_col68[64];
   data_col68[66] <= data_col68[65];
   data_col68[67] <= data_col68[66];
   data_col68[68] <= data_col68[67];

   data_col69[1] <= data[96];
   data_col69[2] <= data_col69[1];
   data_col69[3] <= data_col69[2];
   data_col69[4] <= data_col69[3];
   data_col69[5] <= data_col69[4];
   data_col69[6] <= data_col69[5];
   data_col69[7] <= data_col69[6];
   data_col69[8] <= data_col69[7];
   data_col69[9] <= data_col69[8];
   data_col69[10] <= data_col69[9];
   data_col69[11] <= data_col69[10];
   data_col69[12] <= data_col69[11];
   data_col69[13] <= data_col69[12];
   data_col69[14] <= data_col69[13];
   data_col69[15] <= data_col69[14];
   data_col69[16] <= data_col69[15];
   data_col69[17] <= data_col69[16];
   data_col69[18] <= data_col69[17];
   data_col69[19] <= data_col69[18];
   data_col69[20] <= data_col69[19];
   data_col69[21] <= data_col69[20];
   data_col69[22] <= data_col69[21];
   data_col69[23] <= data_col69[22];
   data_col69[24] <= data_col69[23];
   data_col69[25] <= data_col69[24];
   data_col69[26] <= data_col69[25];
   data_col69[27] <= data_col69[26];
   data_col69[28] <= data_col69[27];
   data_col69[29] <= data_col69[28];
   data_col69[30] <= data_col69[29];
   data_col69[31] <= data_col69[30];
   data_col69[32] <= data_col69[31];
   data_col69[33] <= data_col69[32];
   data_col69[34] <= data_col69[33];
   data_col69[35] <= data_col69[34];
   data_col69[36] <= data_col69[35];
   data_col69[37] <= data_col69[36];
   data_col69[38] <= data_col69[37];
   data_col69[39] <= data_col69[38];
   data_col69[40] <= data_col69[39];
   data_col69[41] <= data_col69[40];
   data_col69[42] <= data_col69[41];
   data_col69[43] <= data_col69[42];
   data_col69[44] <= data_col69[43];
   data_col69[45] <= data_col69[44];
   data_col69[46] <= data_col69[45];
   data_col69[47] <= data_col69[46];
   data_col69[48] <= data_col69[47];
   data_col69[49] <= data_col69[48];
   data_col69[50] <= data_col69[49];
   data_col69[51] <= data_col69[50];
   data_col69[52] <= data_col69[51];
   data_col69[53] <= data_col69[52];
   data_col69[54] <= data_col69[53];
   data_col69[55] <= data_col69[54];
   data_col69[56] <= data_col69[55];
   data_col69[57] <= data_col69[56];
   data_col69[58] <= data_col69[57];
   data_col69[59] <= data_col69[58];
   data_col69[60] <= data_col69[59];
   data_col69[61] <= data_col69[60];
   data_col69[62] <= data_col69[61];
   data_col69[63] <= data_col69[62];
   data_col69[64] <= data_col69[63];
   data_col69[65] <= data_col69[64];
   data_col69[66] <= data_col69[65];
   data_col69[67] <= data_col69[66];
   data_col69[68] <= data_col69[67];
   data_col69[69] <= data_col69[68];

   data_col70[1] <= data[95];
   data_col70[2] <= data_col70[1];
   data_col70[3] <= data_col70[2];
   data_col70[4] <= data_col70[3];
   data_col70[5] <= data_col70[4];
   data_col70[6] <= data_col70[5];
   data_col70[7] <= data_col70[6];
   data_col70[8] <= data_col70[7];
   data_col70[9] <= data_col70[8];
   data_col70[10] <= data_col70[9];
   data_col70[11] <= data_col70[10];
   data_col70[12] <= data_col70[11];
   data_col70[13] <= data_col70[12];
   data_col70[14] <= data_col70[13];
   data_col70[15] <= data_col70[14];
   data_col70[16] <= data_col70[15];
   data_col70[17] <= data_col70[16];
   data_col70[18] <= data_col70[17];
   data_col70[19] <= data_col70[18];
   data_col70[20] <= data_col70[19];
   data_col70[21] <= data_col70[20];
   data_col70[22] <= data_col70[21];
   data_col70[23] <= data_col70[22];
   data_col70[24] <= data_col70[23];
   data_col70[25] <= data_col70[24];
   data_col70[26] <= data_col70[25];
   data_col70[27] <= data_col70[26];
   data_col70[28] <= data_col70[27];
   data_col70[29] <= data_col70[28];
   data_col70[30] <= data_col70[29];
   data_col70[31] <= data_col70[30];
   data_col70[32] <= data_col70[31];
   data_col70[33] <= data_col70[32];
   data_col70[34] <= data_col70[33];
   data_col70[35] <= data_col70[34];
   data_col70[36] <= data_col70[35];
   data_col70[37] <= data_col70[36];
   data_col70[38] <= data_col70[37];
   data_col70[39] <= data_col70[38];
   data_col70[40] <= data_col70[39];
   data_col70[41] <= data_col70[40];
   data_col70[42] <= data_col70[41];
   data_col70[43] <= data_col70[42];
   data_col70[44] <= data_col70[43];
   data_col70[45] <= data_col70[44];
   data_col70[46] <= data_col70[45];
   data_col70[47] <= data_col70[46];
   data_col70[48] <= data_col70[47];
   data_col70[49] <= data_col70[48];
   data_col70[50] <= data_col70[49];
   data_col70[51] <= data_col70[50];
   data_col70[52] <= data_col70[51];
   data_col70[53] <= data_col70[52];
   data_col70[54] <= data_col70[53];
   data_col70[55] <= data_col70[54];
   data_col70[56] <= data_col70[55];
   data_col70[57] <= data_col70[56];
   data_col70[58] <= data_col70[57];
   data_col70[59] <= data_col70[58];
   data_col70[60] <= data_col70[59];
   data_col70[61] <= data_col70[60];
   data_col70[62] <= data_col70[61];
   data_col70[63] <= data_col70[62];
   data_col70[64] <= data_col70[63];
   data_col70[65] <= data_col70[64];
   data_col70[66] <= data_col70[65];
   data_col70[67] <= data_col70[66];
   data_col70[68] <= data_col70[67];
   data_col70[69] <= data_col70[68];
   data_col70[70] <= data_col70[69];

   data_col71[1] <= data[94];
   data_col71[2] <= data_col71[1];
   data_col71[3] <= data_col71[2];
   data_col71[4] <= data_col71[3];
   data_col71[5] <= data_col71[4];
   data_col71[6] <= data_col71[5];
   data_col71[7] <= data_col71[6];
   data_col71[8] <= data_col71[7];
   data_col71[9] <= data_col71[8];
   data_col71[10] <= data_col71[9];
   data_col71[11] <= data_col71[10];
   data_col71[12] <= data_col71[11];
   data_col71[13] <= data_col71[12];
   data_col71[14] <= data_col71[13];
   data_col71[15] <= data_col71[14];
   data_col71[16] <= data_col71[15];
   data_col71[17] <= data_col71[16];
   data_col71[18] <= data_col71[17];
   data_col71[19] <= data_col71[18];
   data_col71[20] <= data_col71[19];
   data_col71[21] <= data_col71[20];
   data_col71[22] <= data_col71[21];
   data_col71[23] <= data_col71[22];
   data_col71[24] <= data_col71[23];
   data_col71[25] <= data_col71[24];
   data_col71[26] <= data_col71[25];
   data_col71[27] <= data_col71[26];
   data_col71[28] <= data_col71[27];
   data_col71[29] <= data_col71[28];
   data_col71[30] <= data_col71[29];
   data_col71[31] <= data_col71[30];
   data_col71[32] <= data_col71[31];
   data_col71[33] <= data_col71[32];
   data_col71[34] <= data_col71[33];
   data_col71[35] <= data_col71[34];
   data_col71[36] <= data_col71[35];
   data_col71[37] <= data_col71[36];
   data_col71[38] <= data_col71[37];
   data_col71[39] <= data_col71[38];
   data_col71[40] <= data_col71[39];
   data_col71[41] <= data_col71[40];
   data_col71[42] <= data_col71[41];
   data_col71[43] <= data_col71[42];
   data_col71[44] <= data_col71[43];
   data_col71[45] <= data_col71[44];
   data_col71[46] <= data_col71[45];
   data_col71[47] <= data_col71[46];
   data_col71[48] <= data_col71[47];
   data_col71[49] <= data_col71[48];
   data_col71[50] <= data_col71[49];
   data_col71[51] <= data_col71[50];
   data_col71[52] <= data_col71[51];
   data_col71[53] <= data_col71[52];
   data_col71[54] <= data_col71[53];
   data_col71[55] <= data_col71[54];
   data_col71[56] <= data_col71[55];
   data_col71[57] <= data_col71[56];
   data_col71[58] <= data_col71[57];
   data_col71[59] <= data_col71[58];
   data_col71[60] <= data_col71[59];
   data_col71[61] <= data_col71[60];
   data_col71[62] <= data_col71[61];
   data_col71[63] <= data_col71[62];
   data_col71[64] <= data_col71[63];
   data_col71[65] <= data_col71[64];
   data_col71[66] <= data_col71[65];
   data_col71[67] <= data_col71[66];
   data_col71[68] <= data_col71[67];
   data_col71[69] <= data_col71[68];
   data_col71[70] <= data_col71[69];
   data_col71[71] <= data_col71[70];

   data_col72[1] <= data[93];
   data_col72[2] <= data_col72[1];
   data_col72[3] <= data_col72[2];
   data_col72[4] <= data_col72[3];
   data_col72[5] <= data_col72[4];
   data_col72[6] <= data_col72[5];
   data_col72[7] <= data_col72[6];
   data_col72[8] <= data_col72[7];
   data_col72[9] <= data_col72[8];
   data_col72[10] <= data_col72[9];
   data_col72[11] <= data_col72[10];
   data_col72[12] <= data_col72[11];
   data_col72[13] <= data_col72[12];
   data_col72[14] <= data_col72[13];
   data_col72[15] <= data_col72[14];
   data_col72[16] <= data_col72[15];
   data_col72[17] <= data_col72[16];
   data_col72[18] <= data_col72[17];
   data_col72[19] <= data_col72[18];
   data_col72[20] <= data_col72[19];
   data_col72[21] <= data_col72[20];
   data_col72[22] <= data_col72[21];
   data_col72[23] <= data_col72[22];
   data_col72[24] <= data_col72[23];
   data_col72[25] <= data_col72[24];
   data_col72[26] <= data_col72[25];
   data_col72[27] <= data_col72[26];
   data_col72[28] <= data_col72[27];
   data_col72[29] <= data_col72[28];
   data_col72[30] <= data_col72[29];
   data_col72[31] <= data_col72[30];
   data_col72[32] <= data_col72[31];
   data_col72[33] <= data_col72[32];
   data_col72[34] <= data_col72[33];
   data_col72[35] <= data_col72[34];
   data_col72[36] <= data_col72[35];
   data_col72[37] <= data_col72[36];
   data_col72[38] <= data_col72[37];
   data_col72[39] <= data_col72[38];
   data_col72[40] <= data_col72[39];
   data_col72[41] <= data_col72[40];
   data_col72[42] <= data_col72[41];
   data_col72[43] <= data_col72[42];
   data_col72[44] <= data_col72[43];
   data_col72[45] <= data_col72[44];
   data_col72[46] <= data_col72[45];
   data_col72[47] <= data_col72[46];
   data_col72[48] <= data_col72[47];
   data_col72[49] <= data_col72[48];
   data_col72[50] <= data_col72[49];
   data_col72[51] <= data_col72[50];
   data_col72[52] <= data_col72[51];
   data_col72[53] <= data_col72[52];
   data_col72[54] <= data_col72[53];
   data_col72[55] <= data_col72[54];
   data_col72[56] <= data_col72[55];
   data_col72[57] <= data_col72[56];
   data_col72[58] <= data_col72[57];
   data_col72[59] <= data_col72[58];
   data_col72[60] <= data_col72[59];
   data_col72[61] <= data_col72[60];
   data_col72[62] <= data_col72[61];
   data_col72[63] <= data_col72[62];
   data_col72[64] <= data_col72[63];
   data_col72[65] <= data_col72[64];
   data_col72[66] <= data_col72[65];
   data_col72[67] <= data_col72[66];
   data_col72[68] <= data_col72[67];
   data_col72[69] <= data_col72[68];
   data_col72[70] <= data_col72[69];
   data_col72[71] <= data_col72[70];
   data_col72[72] <= data_col72[71];

   data_col73[1] <= data[92];
   data_col73[2] <= data_col73[1];
   data_col73[3] <= data_col73[2];
   data_col73[4] <= data_col73[3];
   data_col73[5] <= data_col73[4];
   data_col73[6] <= data_col73[5];
   data_col73[7] <= data_col73[6];
   data_col73[8] <= data_col73[7];
   data_col73[9] <= data_col73[8];
   data_col73[10] <= data_col73[9];
   data_col73[11] <= data_col73[10];
   data_col73[12] <= data_col73[11];
   data_col73[13] <= data_col73[12];
   data_col73[14] <= data_col73[13];
   data_col73[15] <= data_col73[14];
   data_col73[16] <= data_col73[15];
   data_col73[17] <= data_col73[16];
   data_col73[18] <= data_col73[17];
   data_col73[19] <= data_col73[18];
   data_col73[20] <= data_col73[19];
   data_col73[21] <= data_col73[20];
   data_col73[22] <= data_col73[21];
   data_col73[23] <= data_col73[22];
   data_col73[24] <= data_col73[23];
   data_col73[25] <= data_col73[24];
   data_col73[26] <= data_col73[25];
   data_col73[27] <= data_col73[26];
   data_col73[28] <= data_col73[27];
   data_col73[29] <= data_col73[28];
   data_col73[30] <= data_col73[29];
   data_col73[31] <= data_col73[30];
   data_col73[32] <= data_col73[31];
   data_col73[33] <= data_col73[32];
   data_col73[34] <= data_col73[33];
   data_col73[35] <= data_col73[34];
   data_col73[36] <= data_col73[35];
   data_col73[37] <= data_col73[36];
   data_col73[38] <= data_col73[37];
   data_col73[39] <= data_col73[38];
   data_col73[40] <= data_col73[39];
   data_col73[41] <= data_col73[40];
   data_col73[42] <= data_col73[41];
   data_col73[43] <= data_col73[42];
   data_col73[44] <= data_col73[43];
   data_col73[45] <= data_col73[44];
   data_col73[46] <= data_col73[45];
   data_col73[47] <= data_col73[46];
   data_col73[48] <= data_col73[47];
   data_col73[49] <= data_col73[48];
   data_col73[50] <= data_col73[49];
   data_col73[51] <= data_col73[50];
   data_col73[52] <= data_col73[51];
   data_col73[53] <= data_col73[52];
   data_col73[54] <= data_col73[53];
   data_col73[55] <= data_col73[54];
   data_col73[56] <= data_col73[55];
   data_col73[57] <= data_col73[56];
   data_col73[58] <= data_col73[57];
   data_col73[59] <= data_col73[58];
   data_col73[60] <= data_col73[59];
   data_col73[61] <= data_col73[60];
   data_col73[62] <= data_col73[61];
   data_col73[63] <= data_col73[62];
   data_col73[64] <= data_col73[63];
   data_col73[65] <= data_col73[64];
   data_col73[66] <= data_col73[65];
   data_col73[67] <= data_col73[66];
   data_col73[68] <= data_col73[67];
   data_col73[69] <= data_col73[68];
   data_col73[70] <= data_col73[69];
   data_col73[71] <= data_col73[70];
   data_col73[72] <= data_col73[71];
   data_col73[73] <= data_col73[72];

   data_col74[1] <= data[91];
   data_col74[2] <= data_col74[1];
   data_col74[3] <= data_col74[2];
   data_col74[4] <= data_col74[3];
   data_col74[5] <= data_col74[4];
   data_col74[6] <= data_col74[5];
   data_col74[7] <= data_col74[6];
   data_col74[8] <= data_col74[7];
   data_col74[9] <= data_col74[8];
   data_col74[10] <= data_col74[9];
   data_col74[11] <= data_col74[10];
   data_col74[12] <= data_col74[11];
   data_col74[13] <= data_col74[12];
   data_col74[14] <= data_col74[13];
   data_col74[15] <= data_col74[14];
   data_col74[16] <= data_col74[15];
   data_col74[17] <= data_col74[16];
   data_col74[18] <= data_col74[17];
   data_col74[19] <= data_col74[18];
   data_col74[20] <= data_col74[19];
   data_col74[21] <= data_col74[20];
   data_col74[22] <= data_col74[21];
   data_col74[23] <= data_col74[22];
   data_col74[24] <= data_col74[23];
   data_col74[25] <= data_col74[24];
   data_col74[26] <= data_col74[25];
   data_col74[27] <= data_col74[26];
   data_col74[28] <= data_col74[27];
   data_col74[29] <= data_col74[28];
   data_col74[30] <= data_col74[29];
   data_col74[31] <= data_col74[30];
   data_col74[32] <= data_col74[31];
   data_col74[33] <= data_col74[32];
   data_col74[34] <= data_col74[33];
   data_col74[35] <= data_col74[34];
   data_col74[36] <= data_col74[35];
   data_col74[37] <= data_col74[36];
   data_col74[38] <= data_col74[37];
   data_col74[39] <= data_col74[38];
   data_col74[40] <= data_col74[39];
   data_col74[41] <= data_col74[40];
   data_col74[42] <= data_col74[41];
   data_col74[43] <= data_col74[42];
   data_col74[44] <= data_col74[43];
   data_col74[45] <= data_col74[44];
   data_col74[46] <= data_col74[45];
   data_col74[47] <= data_col74[46];
   data_col74[48] <= data_col74[47];
   data_col74[49] <= data_col74[48];
   data_col74[50] <= data_col74[49];
   data_col74[51] <= data_col74[50];
   data_col74[52] <= data_col74[51];
   data_col74[53] <= data_col74[52];
   data_col74[54] <= data_col74[53];
   data_col74[55] <= data_col74[54];
   data_col74[56] <= data_col74[55];
   data_col74[57] <= data_col74[56];
   data_col74[58] <= data_col74[57];
   data_col74[59] <= data_col74[58];
   data_col74[60] <= data_col74[59];
   data_col74[61] <= data_col74[60];
   data_col74[62] <= data_col74[61];
   data_col74[63] <= data_col74[62];
   data_col74[64] <= data_col74[63];
   data_col74[65] <= data_col74[64];
   data_col74[66] <= data_col74[65];
   data_col74[67] <= data_col74[66];
   data_col74[68] <= data_col74[67];
   data_col74[69] <= data_col74[68];
   data_col74[70] <= data_col74[69];
   data_col74[71] <= data_col74[70];
   data_col74[72] <= data_col74[71];
   data_col74[73] <= data_col74[72];
   data_col74[74] <= data_col74[73];

   data_col75[1] <= data[90];
   data_col75[2] <= data_col75[1];
   data_col75[3] <= data_col75[2];
   data_col75[4] <= data_col75[3];
   data_col75[5] <= data_col75[4];
   data_col75[6] <= data_col75[5];
   data_col75[7] <= data_col75[6];
   data_col75[8] <= data_col75[7];
   data_col75[9] <= data_col75[8];
   data_col75[10] <= data_col75[9];
   data_col75[11] <= data_col75[10];
   data_col75[12] <= data_col75[11];
   data_col75[13] <= data_col75[12];
   data_col75[14] <= data_col75[13];
   data_col75[15] <= data_col75[14];
   data_col75[16] <= data_col75[15];
   data_col75[17] <= data_col75[16];
   data_col75[18] <= data_col75[17];
   data_col75[19] <= data_col75[18];
   data_col75[20] <= data_col75[19];
   data_col75[21] <= data_col75[20];
   data_col75[22] <= data_col75[21];
   data_col75[23] <= data_col75[22];
   data_col75[24] <= data_col75[23];
   data_col75[25] <= data_col75[24];
   data_col75[26] <= data_col75[25];
   data_col75[27] <= data_col75[26];
   data_col75[28] <= data_col75[27];
   data_col75[29] <= data_col75[28];
   data_col75[30] <= data_col75[29];
   data_col75[31] <= data_col75[30];
   data_col75[32] <= data_col75[31];
   data_col75[33] <= data_col75[32];
   data_col75[34] <= data_col75[33];
   data_col75[35] <= data_col75[34];
   data_col75[36] <= data_col75[35];
   data_col75[37] <= data_col75[36];
   data_col75[38] <= data_col75[37];
   data_col75[39] <= data_col75[38];
   data_col75[40] <= data_col75[39];
   data_col75[41] <= data_col75[40];
   data_col75[42] <= data_col75[41];
   data_col75[43] <= data_col75[42];
   data_col75[44] <= data_col75[43];
   data_col75[45] <= data_col75[44];
   data_col75[46] <= data_col75[45];
   data_col75[47] <= data_col75[46];
   data_col75[48] <= data_col75[47];
   data_col75[49] <= data_col75[48];
   data_col75[50] <= data_col75[49];
   data_col75[51] <= data_col75[50];
   data_col75[52] <= data_col75[51];
   data_col75[53] <= data_col75[52];
   data_col75[54] <= data_col75[53];
   data_col75[55] <= data_col75[54];
   data_col75[56] <= data_col75[55];
   data_col75[57] <= data_col75[56];
   data_col75[58] <= data_col75[57];
   data_col75[59] <= data_col75[58];
   data_col75[60] <= data_col75[59];
   data_col75[61] <= data_col75[60];
   data_col75[62] <= data_col75[61];
   data_col75[63] <= data_col75[62];
   data_col75[64] <= data_col75[63];
   data_col75[65] <= data_col75[64];
   data_col75[66] <= data_col75[65];
   data_col75[67] <= data_col75[66];
   data_col75[68] <= data_col75[67];
   data_col75[69] <= data_col75[68];
   data_col75[70] <= data_col75[69];
   data_col75[71] <= data_col75[70];
   data_col75[72] <= data_col75[71];
   data_col75[73] <= data_col75[72];
   data_col75[74] <= data_col75[73];
   data_col75[75] <= data_col75[74];

   data_col76[1] <= data[89];
   data_col76[2] <= data_col76[1];
   data_col76[3] <= data_col76[2];
   data_col76[4] <= data_col76[3];
   data_col76[5] <= data_col76[4];
   data_col76[6] <= data_col76[5];
   data_col76[7] <= data_col76[6];
   data_col76[8] <= data_col76[7];
   data_col76[9] <= data_col76[8];
   data_col76[10] <= data_col76[9];
   data_col76[11] <= data_col76[10];
   data_col76[12] <= data_col76[11];
   data_col76[13] <= data_col76[12];
   data_col76[14] <= data_col76[13];
   data_col76[15] <= data_col76[14];
   data_col76[16] <= data_col76[15];
   data_col76[17] <= data_col76[16];
   data_col76[18] <= data_col76[17];
   data_col76[19] <= data_col76[18];
   data_col76[20] <= data_col76[19];
   data_col76[21] <= data_col76[20];
   data_col76[22] <= data_col76[21];
   data_col76[23] <= data_col76[22];
   data_col76[24] <= data_col76[23];
   data_col76[25] <= data_col76[24];
   data_col76[26] <= data_col76[25];
   data_col76[27] <= data_col76[26];
   data_col76[28] <= data_col76[27];
   data_col76[29] <= data_col76[28];
   data_col76[30] <= data_col76[29];
   data_col76[31] <= data_col76[30];
   data_col76[32] <= data_col76[31];
   data_col76[33] <= data_col76[32];
   data_col76[34] <= data_col76[33];
   data_col76[35] <= data_col76[34];
   data_col76[36] <= data_col76[35];
   data_col76[37] <= data_col76[36];
   data_col76[38] <= data_col76[37];
   data_col76[39] <= data_col76[38];
   data_col76[40] <= data_col76[39];
   data_col76[41] <= data_col76[40];
   data_col76[42] <= data_col76[41];
   data_col76[43] <= data_col76[42];
   data_col76[44] <= data_col76[43];
   data_col76[45] <= data_col76[44];
   data_col76[46] <= data_col76[45];
   data_col76[47] <= data_col76[46];
   data_col76[48] <= data_col76[47];
   data_col76[49] <= data_col76[48];
   data_col76[50] <= data_col76[49];
   data_col76[51] <= data_col76[50];
   data_col76[52] <= data_col76[51];
   data_col76[53] <= data_col76[52];
   data_col76[54] <= data_col76[53];
   data_col76[55] <= data_col76[54];
   data_col76[56] <= data_col76[55];
   data_col76[57] <= data_col76[56];
   data_col76[58] <= data_col76[57];
   data_col76[59] <= data_col76[58];
   data_col76[60] <= data_col76[59];
   data_col76[61] <= data_col76[60];
   data_col76[62] <= data_col76[61];
   data_col76[63] <= data_col76[62];
   data_col76[64] <= data_col76[63];
   data_col76[65] <= data_col76[64];
   data_col76[66] <= data_col76[65];
   data_col76[67] <= data_col76[66];
   data_col76[68] <= data_col76[67];
   data_col76[69] <= data_col76[68];
   data_col76[70] <= data_col76[69];
   data_col76[71] <= data_col76[70];
   data_col76[72] <= data_col76[71];
   data_col76[73] <= data_col76[72];
   data_col76[74] <= data_col76[73];
   data_col76[75] <= data_col76[74];
   data_col76[76] <= data_col76[75];

   data_col77[1] <= data[88];
   data_col77[2] <= data_col77[1];
   data_col77[3] <= data_col77[2];
   data_col77[4] <= data_col77[3];
   data_col77[5] <= data_col77[4];
   data_col77[6] <= data_col77[5];
   data_col77[7] <= data_col77[6];
   data_col77[8] <= data_col77[7];
   data_col77[9] <= data_col77[8];
   data_col77[10] <= data_col77[9];
   data_col77[11] <= data_col77[10];
   data_col77[12] <= data_col77[11];
   data_col77[13] <= data_col77[12];
   data_col77[14] <= data_col77[13];
   data_col77[15] <= data_col77[14];
   data_col77[16] <= data_col77[15];
   data_col77[17] <= data_col77[16];
   data_col77[18] <= data_col77[17];
   data_col77[19] <= data_col77[18];
   data_col77[20] <= data_col77[19];
   data_col77[21] <= data_col77[20];
   data_col77[22] <= data_col77[21];
   data_col77[23] <= data_col77[22];
   data_col77[24] <= data_col77[23];
   data_col77[25] <= data_col77[24];
   data_col77[26] <= data_col77[25];
   data_col77[27] <= data_col77[26];
   data_col77[28] <= data_col77[27];
   data_col77[29] <= data_col77[28];
   data_col77[30] <= data_col77[29];
   data_col77[31] <= data_col77[30];
   data_col77[32] <= data_col77[31];
   data_col77[33] <= data_col77[32];
   data_col77[34] <= data_col77[33];
   data_col77[35] <= data_col77[34];
   data_col77[36] <= data_col77[35];
   data_col77[37] <= data_col77[36];
   data_col77[38] <= data_col77[37];
   data_col77[39] <= data_col77[38];
   data_col77[40] <= data_col77[39];
   data_col77[41] <= data_col77[40];
   data_col77[42] <= data_col77[41];
   data_col77[43] <= data_col77[42];
   data_col77[44] <= data_col77[43];
   data_col77[45] <= data_col77[44];
   data_col77[46] <= data_col77[45];
   data_col77[47] <= data_col77[46];
   data_col77[48] <= data_col77[47];
   data_col77[49] <= data_col77[48];
   data_col77[50] <= data_col77[49];
   data_col77[51] <= data_col77[50];
   data_col77[52] <= data_col77[51];
   data_col77[53] <= data_col77[52];
   data_col77[54] <= data_col77[53];
   data_col77[55] <= data_col77[54];
   data_col77[56] <= data_col77[55];
   data_col77[57] <= data_col77[56];
   data_col77[58] <= data_col77[57];
   data_col77[59] <= data_col77[58];
   data_col77[60] <= data_col77[59];
   data_col77[61] <= data_col77[60];
   data_col77[62] <= data_col77[61];
   data_col77[63] <= data_col77[62];
   data_col77[64] <= data_col77[63];
   data_col77[65] <= data_col77[64];
   data_col77[66] <= data_col77[65];
   data_col77[67] <= data_col77[66];
   data_col77[68] <= data_col77[67];
   data_col77[69] <= data_col77[68];
   data_col77[70] <= data_col77[69];
   data_col77[71] <= data_col77[70];
   data_col77[72] <= data_col77[71];
   data_col77[73] <= data_col77[72];
   data_col77[74] <= data_col77[73];
   data_col77[75] <= data_col77[74];
   data_col77[76] <= data_col77[75];
   data_col77[77] <= data_col77[76];

   data_col78[1] <= data[87];
   data_col78[2] <= data_col78[1];
   data_col78[3] <= data_col78[2];
   data_col78[4] <= data_col78[3];
   data_col78[5] <= data_col78[4];
   data_col78[6] <= data_col78[5];
   data_col78[7] <= data_col78[6];
   data_col78[8] <= data_col78[7];
   data_col78[9] <= data_col78[8];
   data_col78[10] <= data_col78[9];
   data_col78[11] <= data_col78[10];
   data_col78[12] <= data_col78[11];
   data_col78[13] <= data_col78[12];
   data_col78[14] <= data_col78[13];
   data_col78[15] <= data_col78[14];
   data_col78[16] <= data_col78[15];
   data_col78[17] <= data_col78[16];
   data_col78[18] <= data_col78[17];
   data_col78[19] <= data_col78[18];
   data_col78[20] <= data_col78[19];
   data_col78[21] <= data_col78[20];
   data_col78[22] <= data_col78[21];
   data_col78[23] <= data_col78[22];
   data_col78[24] <= data_col78[23];
   data_col78[25] <= data_col78[24];
   data_col78[26] <= data_col78[25];
   data_col78[27] <= data_col78[26];
   data_col78[28] <= data_col78[27];
   data_col78[29] <= data_col78[28];
   data_col78[30] <= data_col78[29];
   data_col78[31] <= data_col78[30];
   data_col78[32] <= data_col78[31];
   data_col78[33] <= data_col78[32];
   data_col78[34] <= data_col78[33];
   data_col78[35] <= data_col78[34];
   data_col78[36] <= data_col78[35];
   data_col78[37] <= data_col78[36];
   data_col78[38] <= data_col78[37];
   data_col78[39] <= data_col78[38];
   data_col78[40] <= data_col78[39];
   data_col78[41] <= data_col78[40];
   data_col78[42] <= data_col78[41];
   data_col78[43] <= data_col78[42];
   data_col78[44] <= data_col78[43];
   data_col78[45] <= data_col78[44];
   data_col78[46] <= data_col78[45];
   data_col78[47] <= data_col78[46];
   data_col78[48] <= data_col78[47];
   data_col78[49] <= data_col78[48];
   data_col78[50] <= data_col78[49];
   data_col78[51] <= data_col78[50];
   data_col78[52] <= data_col78[51];
   data_col78[53] <= data_col78[52];
   data_col78[54] <= data_col78[53];
   data_col78[55] <= data_col78[54];
   data_col78[56] <= data_col78[55];
   data_col78[57] <= data_col78[56];
   data_col78[58] <= data_col78[57];
   data_col78[59] <= data_col78[58];
   data_col78[60] <= data_col78[59];
   data_col78[61] <= data_col78[60];
   data_col78[62] <= data_col78[61];
   data_col78[63] <= data_col78[62];
   data_col78[64] <= data_col78[63];
   data_col78[65] <= data_col78[64];
   data_col78[66] <= data_col78[65];
   data_col78[67] <= data_col78[66];
   data_col78[68] <= data_col78[67];
   data_col78[69] <= data_col78[68];
   data_col78[70] <= data_col78[69];
   data_col78[71] <= data_col78[70];
   data_col78[72] <= data_col78[71];
   data_col78[73] <= data_col78[72];
   data_col78[74] <= data_col78[73];
   data_col78[75] <= data_col78[74];
   data_col78[76] <= data_col78[75];
   data_col78[77] <= data_col78[76];
   data_col78[78] <= data_col78[77];

   data_col79[1] <= data[86];
   data_col79[2] <= data_col79[1];
   data_col79[3] <= data_col79[2];
   data_col79[4] <= data_col79[3];
   data_col79[5] <= data_col79[4];
   data_col79[6] <= data_col79[5];
   data_col79[7] <= data_col79[6];
   data_col79[8] <= data_col79[7];
   data_col79[9] <= data_col79[8];
   data_col79[10] <= data_col79[9];
   data_col79[11] <= data_col79[10];
   data_col79[12] <= data_col79[11];
   data_col79[13] <= data_col79[12];
   data_col79[14] <= data_col79[13];
   data_col79[15] <= data_col79[14];
   data_col79[16] <= data_col79[15];
   data_col79[17] <= data_col79[16];
   data_col79[18] <= data_col79[17];
   data_col79[19] <= data_col79[18];
   data_col79[20] <= data_col79[19];
   data_col79[21] <= data_col79[20];
   data_col79[22] <= data_col79[21];
   data_col79[23] <= data_col79[22];
   data_col79[24] <= data_col79[23];
   data_col79[25] <= data_col79[24];
   data_col79[26] <= data_col79[25];
   data_col79[27] <= data_col79[26];
   data_col79[28] <= data_col79[27];
   data_col79[29] <= data_col79[28];
   data_col79[30] <= data_col79[29];
   data_col79[31] <= data_col79[30];
   data_col79[32] <= data_col79[31];
   data_col79[33] <= data_col79[32];
   data_col79[34] <= data_col79[33];
   data_col79[35] <= data_col79[34];
   data_col79[36] <= data_col79[35];
   data_col79[37] <= data_col79[36];
   data_col79[38] <= data_col79[37];
   data_col79[39] <= data_col79[38];
   data_col79[40] <= data_col79[39];
   data_col79[41] <= data_col79[40];
   data_col79[42] <= data_col79[41];
   data_col79[43] <= data_col79[42];
   data_col79[44] <= data_col79[43];
   data_col79[45] <= data_col79[44];
   data_col79[46] <= data_col79[45];
   data_col79[47] <= data_col79[46];
   data_col79[48] <= data_col79[47];
   data_col79[49] <= data_col79[48];
   data_col79[50] <= data_col79[49];
   data_col79[51] <= data_col79[50];
   data_col79[52] <= data_col79[51];
   data_col79[53] <= data_col79[52];
   data_col79[54] <= data_col79[53];
   data_col79[55] <= data_col79[54];
   data_col79[56] <= data_col79[55];
   data_col79[57] <= data_col79[56];
   data_col79[58] <= data_col79[57];
   data_col79[59] <= data_col79[58];
   data_col79[60] <= data_col79[59];
   data_col79[61] <= data_col79[60];
   data_col79[62] <= data_col79[61];
   data_col79[63] <= data_col79[62];
   data_col79[64] <= data_col79[63];
   data_col79[65] <= data_col79[64];
   data_col79[66] <= data_col79[65];
   data_col79[67] <= data_col79[66];
   data_col79[68] <= data_col79[67];
   data_col79[69] <= data_col79[68];
   data_col79[70] <= data_col79[69];
   data_col79[71] <= data_col79[70];
   data_col79[72] <= data_col79[71];
   data_col79[73] <= data_col79[72];
   data_col79[74] <= data_col79[73];
   data_col79[75] <= data_col79[74];
   data_col79[76] <= data_col79[75];
   data_col79[77] <= data_col79[76];
   data_col79[78] <= data_col79[77];
   data_col79[79] <= data_col79[78];

   data_col80[1] <= data[85];
   data_col80[2] <= data_col80[1];
   data_col80[3] <= data_col80[2];
   data_col80[4] <= data_col80[3];
   data_col80[5] <= data_col80[4];
   data_col80[6] <= data_col80[5];
   data_col80[7] <= data_col80[6];
   data_col80[8] <= data_col80[7];
   data_col80[9] <= data_col80[8];
   data_col80[10] <= data_col80[9];
   data_col80[11] <= data_col80[10];
   data_col80[12] <= data_col80[11];
   data_col80[13] <= data_col80[12];
   data_col80[14] <= data_col80[13];
   data_col80[15] <= data_col80[14];
   data_col80[16] <= data_col80[15];
   data_col80[17] <= data_col80[16];
   data_col80[18] <= data_col80[17];
   data_col80[19] <= data_col80[18];
   data_col80[20] <= data_col80[19];
   data_col80[21] <= data_col80[20];
   data_col80[22] <= data_col80[21];
   data_col80[23] <= data_col80[22];
   data_col80[24] <= data_col80[23];
   data_col80[25] <= data_col80[24];
   data_col80[26] <= data_col80[25];
   data_col80[27] <= data_col80[26];
   data_col80[28] <= data_col80[27];
   data_col80[29] <= data_col80[28];
   data_col80[30] <= data_col80[29];
   data_col80[31] <= data_col80[30];
   data_col80[32] <= data_col80[31];
   data_col80[33] <= data_col80[32];
   data_col80[34] <= data_col80[33];
   data_col80[35] <= data_col80[34];
   data_col80[36] <= data_col80[35];
   data_col80[37] <= data_col80[36];
   data_col80[38] <= data_col80[37];
   data_col80[39] <= data_col80[38];
   data_col80[40] <= data_col80[39];
   data_col80[41] <= data_col80[40];
   data_col80[42] <= data_col80[41];
   data_col80[43] <= data_col80[42];
   data_col80[44] <= data_col80[43];
   data_col80[45] <= data_col80[44];
   data_col80[46] <= data_col80[45];
   data_col80[47] <= data_col80[46];
   data_col80[48] <= data_col80[47];
   data_col80[49] <= data_col80[48];
   data_col80[50] <= data_col80[49];
   data_col80[51] <= data_col80[50];
   data_col80[52] <= data_col80[51];
   data_col80[53] <= data_col80[52];
   data_col80[54] <= data_col80[53];
   data_col80[55] <= data_col80[54];
   data_col80[56] <= data_col80[55];
   data_col80[57] <= data_col80[56];
   data_col80[58] <= data_col80[57];
   data_col80[59] <= data_col80[58];
   data_col80[60] <= data_col80[59];
   data_col80[61] <= data_col80[60];
   data_col80[62] <= data_col80[61];
   data_col80[63] <= data_col80[62];
   data_col80[64] <= data_col80[63];
   data_col80[65] <= data_col80[64];
   data_col80[66] <= data_col80[65];
   data_col80[67] <= data_col80[66];
   data_col80[68] <= data_col80[67];
   data_col80[69] <= data_col80[68];
   data_col80[70] <= data_col80[69];
   data_col80[71] <= data_col80[70];
   data_col80[72] <= data_col80[71];
   data_col80[73] <= data_col80[72];
   data_col80[74] <= data_col80[73];
   data_col80[75] <= data_col80[74];
   data_col80[76] <= data_col80[75];
   data_col80[77] <= data_col80[76];
   data_col80[78] <= data_col80[77];
   data_col80[79] <= data_col80[78];
   data_col80[80] <= data_col80[79];

   data_col81[1] <= data[84];
   data_col81[2] <= data_col81[1];
   data_col81[3] <= data_col81[2];
   data_col81[4] <= data_col81[3];
   data_col81[5] <= data_col81[4];
   data_col81[6] <= data_col81[5];
   data_col81[7] <= data_col81[6];
   data_col81[8] <= data_col81[7];
   data_col81[9] <= data_col81[8];
   data_col81[10] <= data_col81[9];
   data_col81[11] <= data_col81[10];
   data_col81[12] <= data_col81[11];
   data_col81[13] <= data_col81[12];
   data_col81[14] <= data_col81[13];
   data_col81[15] <= data_col81[14];
   data_col81[16] <= data_col81[15];
   data_col81[17] <= data_col81[16];
   data_col81[18] <= data_col81[17];
   data_col81[19] <= data_col81[18];
   data_col81[20] <= data_col81[19];
   data_col81[21] <= data_col81[20];
   data_col81[22] <= data_col81[21];
   data_col81[23] <= data_col81[22];
   data_col81[24] <= data_col81[23];
   data_col81[25] <= data_col81[24];
   data_col81[26] <= data_col81[25];
   data_col81[27] <= data_col81[26];
   data_col81[28] <= data_col81[27];
   data_col81[29] <= data_col81[28];
   data_col81[30] <= data_col81[29];
   data_col81[31] <= data_col81[30];
   data_col81[32] <= data_col81[31];
   data_col81[33] <= data_col81[32];
   data_col81[34] <= data_col81[33];
   data_col81[35] <= data_col81[34];
   data_col81[36] <= data_col81[35];
   data_col81[37] <= data_col81[36];
   data_col81[38] <= data_col81[37];
   data_col81[39] <= data_col81[38];
   data_col81[40] <= data_col81[39];
   data_col81[41] <= data_col81[40];
   data_col81[42] <= data_col81[41];
   data_col81[43] <= data_col81[42];
   data_col81[44] <= data_col81[43];
   data_col81[45] <= data_col81[44];
   data_col81[46] <= data_col81[45];
   data_col81[47] <= data_col81[46];
   data_col81[48] <= data_col81[47];
   data_col81[49] <= data_col81[48];
   data_col81[50] <= data_col81[49];
   data_col81[51] <= data_col81[50];
   data_col81[52] <= data_col81[51];
   data_col81[53] <= data_col81[52];
   data_col81[54] <= data_col81[53];
   data_col81[55] <= data_col81[54];
   data_col81[56] <= data_col81[55];
   data_col81[57] <= data_col81[56];
   data_col81[58] <= data_col81[57];
   data_col81[59] <= data_col81[58];
   data_col81[60] <= data_col81[59];
   data_col81[61] <= data_col81[60];
   data_col81[62] <= data_col81[61];
   data_col81[63] <= data_col81[62];
   data_col81[64] <= data_col81[63];
   data_col81[65] <= data_col81[64];
   data_col81[66] <= data_col81[65];
   data_col81[67] <= data_col81[66];
   data_col81[68] <= data_col81[67];
   data_col81[69] <= data_col81[68];
   data_col81[70] <= data_col81[69];
   data_col81[71] <= data_col81[70];
   data_col81[72] <= data_col81[71];
   data_col81[73] <= data_col81[72];
   data_col81[74] <= data_col81[73];
   data_col81[75] <= data_col81[74];
   data_col81[76] <= data_col81[75];
   data_col81[77] <= data_col81[76];
   data_col81[78] <= data_col81[77];
   data_col81[79] <= data_col81[78];
   data_col81[80] <= data_col81[79];
   data_col81[81] <= data_col81[80];

   data_col82[1] <= data[83];
   data_col82[2] <= data_col82[1];
   data_col82[3] <= data_col82[2];
   data_col82[4] <= data_col82[3];
   data_col82[5] <= data_col82[4];
   data_col82[6] <= data_col82[5];
   data_col82[7] <= data_col82[6];
   data_col82[8] <= data_col82[7];
   data_col82[9] <= data_col82[8];
   data_col82[10] <= data_col82[9];
   data_col82[11] <= data_col82[10];
   data_col82[12] <= data_col82[11];
   data_col82[13] <= data_col82[12];
   data_col82[14] <= data_col82[13];
   data_col82[15] <= data_col82[14];
   data_col82[16] <= data_col82[15];
   data_col82[17] <= data_col82[16];
   data_col82[18] <= data_col82[17];
   data_col82[19] <= data_col82[18];
   data_col82[20] <= data_col82[19];
   data_col82[21] <= data_col82[20];
   data_col82[22] <= data_col82[21];
   data_col82[23] <= data_col82[22];
   data_col82[24] <= data_col82[23];
   data_col82[25] <= data_col82[24];
   data_col82[26] <= data_col82[25];
   data_col82[27] <= data_col82[26];
   data_col82[28] <= data_col82[27];
   data_col82[29] <= data_col82[28];
   data_col82[30] <= data_col82[29];
   data_col82[31] <= data_col82[30];
   data_col82[32] <= data_col82[31];
   data_col82[33] <= data_col82[32];
   data_col82[34] <= data_col82[33];
   data_col82[35] <= data_col82[34];
   data_col82[36] <= data_col82[35];
   data_col82[37] <= data_col82[36];
   data_col82[38] <= data_col82[37];
   data_col82[39] <= data_col82[38];
   data_col82[40] <= data_col82[39];
   data_col82[41] <= data_col82[40];
   data_col82[42] <= data_col82[41];
   data_col82[43] <= data_col82[42];
   data_col82[44] <= data_col82[43];
   data_col82[45] <= data_col82[44];
   data_col82[46] <= data_col82[45];
   data_col82[47] <= data_col82[46];
   data_col82[48] <= data_col82[47];
   data_col82[49] <= data_col82[48];
   data_col82[50] <= data_col82[49];
   data_col82[51] <= data_col82[50];
   data_col82[52] <= data_col82[51];
   data_col82[53] <= data_col82[52];
   data_col82[54] <= data_col82[53];
   data_col82[55] <= data_col82[54];
   data_col82[56] <= data_col82[55];
   data_col82[57] <= data_col82[56];
   data_col82[58] <= data_col82[57];
   data_col82[59] <= data_col82[58];
   data_col82[60] <= data_col82[59];
   data_col82[61] <= data_col82[60];
   data_col82[62] <= data_col82[61];
   data_col82[63] <= data_col82[62];
   data_col82[64] <= data_col82[63];
   data_col82[65] <= data_col82[64];
   data_col82[66] <= data_col82[65];
   data_col82[67] <= data_col82[66];
   data_col82[68] <= data_col82[67];
   data_col82[69] <= data_col82[68];
   data_col82[70] <= data_col82[69];
   data_col82[71] <= data_col82[70];
   data_col82[72] <= data_col82[71];
   data_col82[73] <= data_col82[72];
   data_col82[74] <= data_col82[73];
   data_col82[75] <= data_col82[74];
   data_col82[76] <= data_col82[75];
   data_col82[77] <= data_col82[76];
   data_col82[78] <= data_col82[77];
   data_col82[79] <= data_col82[78];
   data_col82[80] <= data_col82[79];
   data_col82[81] <= data_col82[80];
   data_col82[82] <= data_col82[81];

   data_col83[1] <= data[82];
   data_col83[2] <= data_col83[1];
   data_col83[3] <= data_col83[2];
   data_col83[4] <= data_col83[3];
   data_col83[5] <= data_col83[4];
   data_col83[6] <= data_col83[5];
   data_col83[7] <= data_col83[6];
   data_col83[8] <= data_col83[7];
   data_col83[9] <= data_col83[8];
   data_col83[10] <= data_col83[9];
   data_col83[11] <= data_col83[10];
   data_col83[12] <= data_col83[11];
   data_col83[13] <= data_col83[12];
   data_col83[14] <= data_col83[13];
   data_col83[15] <= data_col83[14];
   data_col83[16] <= data_col83[15];
   data_col83[17] <= data_col83[16];
   data_col83[18] <= data_col83[17];
   data_col83[19] <= data_col83[18];
   data_col83[20] <= data_col83[19];
   data_col83[21] <= data_col83[20];
   data_col83[22] <= data_col83[21];
   data_col83[23] <= data_col83[22];
   data_col83[24] <= data_col83[23];
   data_col83[25] <= data_col83[24];
   data_col83[26] <= data_col83[25];
   data_col83[27] <= data_col83[26];
   data_col83[28] <= data_col83[27];
   data_col83[29] <= data_col83[28];
   data_col83[30] <= data_col83[29];
   data_col83[31] <= data_col83[30];
   data_col83[32] <= data_col83[31];
   data_col83[33] <= data_col83[32];
   data_col83[34] <= data_col83[33];
   data_col83[35] <= data_col83[34];
   data_col83[36] <= data_col83[35];
   data_col83[37] <= data_col83[36];
   data_col83[38] <= data_col83[37];
   data_col83[39] <= data_col83[38];
   data_col83[40] <= data_col83[39];
   data_col83[41] <= data_col83[40];
   data_col83[42] <= data_col83[41];
   data_col83[43] <= data_col83[42];
   data_col83[44] <= data_col83[43];
   data_col83[45] <= data_col83[44];
   data_col83[46] <= data_col83[45];
   data_col83[47] <= data_col83[46];
   data_col83[48] <= data_col83[47];
   data_col83[49] <= data_col83[48];
   data_col83[50] <= data_col83[49];
   data_col83[51] <= data_col83[50];
   data_col83[52] <= data_col83[51];
   data_col83[53] <= data_col83[52];
   data_col83[54] <= data_col83[53];
   data_col83[55] <= data_col83[54];
   data_col83[56] <= data_col83[55];
   data_col83[57] <= data_col83[56];
   data_col83[58] <= data_col83[57];
   data_col83[59] <= data_col83[58];
   data_col83[60] <= data_col83[59];
   data_col83[61] <= data_col83[60];
   data_col83[62] <= data_col83[61];
   data_col83[63] <= data_col83[62];
   data_col83[64] <= data_col83[63];
   data_col83[65] <= data_col83[64];
   data_col83[66] <= data_col83[65];
   data_col83[67] <= data_col83[66];
   data_col83[68] <= data_col83[67];
   data_col83[69] <= data_col83[68];
   data_col83[70] <= data_col83[69];
   data_col83[71] <= data_col83[70];
   data_col83[72] <= data_col83[71];
   data_col83[73] <= data_col83[72];
   data_col83[74] <= data_col83[73];
   data_col83[75] <= data_col83[74];
   data_col83[76] <= data_col83[75];
   data_col83[77] <= data_col83[76];
   data_col83[78] <= data_col83[77];
   data_col83[79] <= data_col83[78];
   data_col83[80] <= data_col83[79];
   data_col83[81] <= data_col83[80];
   data_col83[82] <= data_col83[81];
   data_col83[83] <= data_col83[82];

   data_col84[1] <= data[81];
   data_col84[2] <= data_col84[1];
   data_col84[3] <= data_col84[2];
   data_col84[4] <= data_col84[3];
   data_col84[5] <= data_col84[4];
   data_col84[6] <= data_col84[5];
   data_col84[7] <= data_col84[6];
   data_col84[8] <= data_col84[7];
   data_col84[9] <= data_col84[8];
   data_col84[10] <= data_col84[9];
   data_col84[11] <= data_col84[10];
   data_col84[12] <= data_col84[11];
   data_col84[13] <= data_col84[12];
   data_col84[14] <= data_col84[13];
   data_col84[15] <= data_col84[14];
   data_col84[16] <= data_col84[15];
   data_col84[17] <= data_col84[16];
   data_col84[18] <= data_col84[17];
   data_col84[19] <= data_col84[18];
   data_col84[20] <= data_col84[19];
   data_col84[21] <= data_col84[20];
   data_col84[22] <= data_col84[21];
   data_col84[23] <= data_col84[22];
   data_col84[24] <= data_col84[23];
   data_col84[25] <= data_col84[24];
   data_col84[26] <= data_col84[25];
   data_col84[27] <= data_col84[26];
   data_col84[28] <= data_col84[27];
   data_col84[29] <= data_col84[28];
   data_col84[30] <= data_col84[29];
   data_col84[31] <= data_col84[30];
   data_col84[32] <= data_col84[31];
   data_col84[33] <= data_col84[32];
   data_col84[34] <= data_col84[33];
   data_col84[35] <= data_col84[34];
   data_col84[36] <= data_col84[35];
   data_col84[37] <= data_col84[36];
   data_col84[38] <= data_col84[37];
   data_col84[39] <= data_col84[38];
   data_col84[40] <= data_col84[39];
   data_col84[41] <= data_col84[40];
   data_col84[42] <= data_col84[41];
   data_col84[43] <= data_col84[42];
   data_col84[44] <= data_col84[43];
   data_col84[45] <= data_col84[44];
   data_col84[46] <= data_col84[45];
   data_col84[47] <= data_col84[46];
   data_col84[48] <= data_col84[47];
   data_col84[49] <= data_col84[48];
   data_col84[50] <= data_col84[49];
   data_col84[51] <= data_col84[50];
   data_col84[52] <= data_col84[51];
   data_col84[53] <= data_col84[52];
   data_col84[54] <= data_col84[53];
   data_col84[55] <= data_col84[54];
   data_col84[56] <= data_col84[55];
   data_col84[57] <= data_col84[56];
   data_col84[58] <= data_col84[57];
   data_col84[59] <= data_col84[58];
   data_col84[60] <= data_col84[59];
   data_col84[61] <= data_col84[60];
   data_col84[62] <= data_col84[61];
   data_col84[63] <= data_col84[62];
   data_col84[64] <= data_col84[63];
   data_col84[65] <= data_col84[64];
   data_col84[66] <= data_col84[65];
   data_col84[67] <= data_col84[66];
   data_col84[68] <= data_col84[67];
   data_col84[69] <= data_col84[68];
   data_col84[70] <= data_col84[69];
   data_col84[71] <= data_col84[70];
   data_col84[72] <= data_col84[71];
   data_col84[73] <= data_col84[72];
   data_col84[74] <= data_col84[73];
   data_col84[75] <= data_col84[74];
   data_col84[76] <= data_col84[75];
   data_col84[77] <= data_col84[76];
   data_col84[78] <= data_col84[77];
   data_col84[79] <= data_col84[78];
   data_col84[80] <= data_col84[79];
   data_col84[81] <= data_col84[80];
   data_col84[82] <= data_col84[81];
   data_col84[83] <= data_col84[82];
   data_col84[84] <= data_col84[83];

   data_col85[1] <= data[80];
   data_col85[2] <= data_col85[1];
   data_col85[3] <= data_col85[2];
   data_col85[4] <= data_col85[3];
   data_col85[5] <= data_col85[4];
   data_col85[6] <= data_col85[5];
   data_col85[7] <= data_col85[6];
   data_col85[8] <= data_col85[7];
   data_col85[9] <= data_col85[8];
   data_col85[10] <= data_col85[9];
   data_col85[11] <= data_col85[10];
   data_col85[12] <= data_col85[11];
   data_col85[13] <= data_col85[12];
   data_col85[14] <= data_col85[13];
   data_col85[15] <= data_col85[14];
   data_col85[16] <= data_col85[15];
   data_col85[17] <= data_col85[16];
   data_col85[18] <= data_col85[17];
   data_col85[19] <= data_col85[18];
   data_col85[20] <= data_col85[19];
   data_col85[21] <= data_col85[20];
   data_col85[22] <= data_col85[21];
   data_col85[23] <= data_col85[22];
   data_col85[24] <= data_col85[23];
   data_col85[25] <= data_col85[24];
   data_col85[26] <= data_col85[25];
   data_col85[27] <= data_col85[26];
   data_col85[28] <= data_col85[27];
   data_col85[29] <= data_col85[28];
   data_col85[30] <= data_col85[29];
   data_col85[31] <= data_col85[30];
   data_col85[32] <= data_col85[31];
   data_col85[33] <= data_col85[32];
   data_col85[34] <= data_col85[33];
   data_col85[35] <= data_col85[34];
   data_col85[36] <= data_col85[35];
   data_col85[37] <= data_col85[36];
   data_col85[38] <= data_col85[37];
   data_col85[39] <= data_col85[38];
   data_col85[40] <= data_col85[39];
   data_col85[41] <= data_col85[40];
   data_col85[42] <= data_col85[41];
   data_col85[43] <= data_col85[42];
   data_col85[44] <= data_col85[43];
   data_col85[45] <= data_col85[44];
   data_col85[46] <= data_col85[45];
   data_col85[47] <= data_col85[46];
   data_col85[48] <= data_col85[47];
   data_col85[49] <= data_col85[48];
   data_col85[50] <= data_col85[49];
   data_col85[51] <= data_col85[50];
   data_col85[52] <= data_col85[51];
   data_col85[53] <= data_col85[52];
   data_col85[54] <= data_col85[53];
   data_col85[55] <= data_col85[54];
   data_col85[56] <= data_col85[55];
   data_col85[57] <= data_col85[56];
   data_col85[58] <= data_col85[57];
   data_col85[59] <= data_col85[58];
   data_col85[60] <= data_col85[59];
   data_col85[61] <= data_col85[60];
   data_col85[62] <= data_col85[61];
   data_col85[63] <= data_col85[62];
   data_col85[64] <= data_col85[63];
   data_col85[65] <= data_col85[64];
   data_col85[66] <= data_col85[65];
   data_col85[67] <= data_col85[66];
   data_col85[68] <= data_col85[67];
   data_col85[69] <= data_col85[68];
   data_col85[70] <= data_col85[69];
   data_col85[71] <= data_col85[70];
   data_col85[72] <= data_col85[71];
   data_col85[73] <= data_col85[72];
   data_col85[74] <= data_col85[73];
   data_col85[75] <= data_col85[74];
   data_col85[76] <= data_col85[75];
   data_col85[77] <= data_col85[76];
   data_col85[78] <= data_col85[77];
   data_col85[79] <= data_col85[78];
   data_col85[80] <= data_col85[79];
   data_col85[81] <= data_col85[80];
   data_col85[82] <= data_col85[81];
   data_col85[83] <= data_col85[82];
   data_col85[84] <= data_col85[83];
   data_col85[85] <= data_col85[84];

   data_col86[1] <= data[79];
   data_col86[2] <= data_col86[1];
   data_col86[3] <= data_col86[2];
   data_col86[4] <= data_col86[3];
   data_col86[5] <= data_col86[4];
   data_col86[6] <= data_col86[5];
   data_col86[7] <= data_col86[6];
   data_col86[8] <= data_col86[7];
   data_col86[9] <= data_col86[8];
   data_col86[10] <= data_col86[9];
   data_col86[11] <= data_col86[10];
   data_col86[12] <= data_col86[11];
   data_col86[13] <= data_col86[12];
   data_col86[14] <= data_col86[13];
   data_col86[15] <= data_col86[14];
   data_col86[16] <= data_col86[15];
   data_col86[17] <= data_col86[16];
   data_col86[18] <= data_col86[17];
   data_col86[19] <= data_col86[18];
   data_col86[20] <= data_col86[19];
   data_col86[21] <= data_col86[20];
   data_col86[22] <= data_col86[21];
   data_col86[23] <= data_col86[22];
   data_col86[24] <= data_col86[23];
   data_col86[25] <= data_col86[24];
   data_col86[26] <= data_col86[25];
   data_col86[27] <= data_col86[26];
   data_col86[28] <= data_col86[27];
   data_col86[29] <= data_col86[28];
   data_col86[30] <= data_col86[29];
   data_col86[31] <= data_col86[30];
   data_col86[32] <= data_col86[31];
   data_col86[33] <= data_col86[32];
   data_col86[34] <= data_col86[33];
   data_col86[35] <= data_col86[34];
   data_col86[36] <= data_col86[35];
   data_col86[37] <= data_col86[36];
   data_col86[38] <= data_col86[37];
   data_col86[39] <= data_col86[38];
   data_col86[40] <= data_col86[39];
   data_col86[41] <= data_col86[40];
   data_col86[42] <= data_col86[41];
   data_col86[43] <= data_col86[42];
   data_col86[44] <= data_col86[43];
   data_col86[45] <= data_col86[44];
   data_col86[46] <= data_col86[45];
   data_col86[47] <= data_col86[46];
   data_col86[48] <= data_col86[47];
   data_col86[49] <= data_col86[48];
   data_col86[50] <= data_col86[49];
   data_col86[51] <= data_col86[50];
   data_col86[52] <= data_col86[51];
   data_col86[53] <= data_col86[52];
   data_col86[54] <= data_col86[53];
   data_col86[55] <= data_col86[54];
   data_col86[56] <= data_col86[55];
   data_col86[57] <= data_col86[56];
   data_col86[58] <= data_col86[57];
   data_col86[59] <= data_col86[58];
   data_col86[60] <= data_col86[59];
   data_col86[61] <= data_col86[60];
   data_col86[62] <= data_col86[61];
   data_col86[63] <= data_col86[62];
   data_col86[64] <= data_col86[63];
   data_col86[65] <= data_col86[64];
   data_col86[66] <= data_col86[65];
   data_col86[67] <= data_col86[66];
   data_col86[68] <= data_col86[67];
   data_col86[69] <= data_col86[68];
   data_col86[70] <= data_col86[69];
   data_col86[71] <= data_col86[70];
   data_col86[72] <= data_col86[71];
   data_col86[73] <= data_col86[72];
   data_col86[74] <= data_col86[73];
   data_col86[75] <= data_col86[74];
   data_col86[76] <= data_col86[75];
   data_col86[77] <= data_col86[76];
   data_col86[78] <= data_col86[77];
   data_col86[79] <= data_col86[78];
   data_col86[80] <= data_col86[79];
   data_col86[81] <= data_col86[80];
   data_col86[82] <= data_col86[81];
   data_col86[83] <= data_col86[82];
   data_col86[84] <= data_col86[83];
   data_col86[85] <= data_col86[84];
   data_col86[86] <= data_col86[85];

   data_col87[1] <= data[78];
   data_col87[2] <= data_col87[1];
   data_col87[3] <= data_col87[2];
   data_col87[4] <= data_col87[3];
   data_col87[5] <= data_col87[4];
   data_col87[6] <= data_col87[5];
   data_col87[7] <= data_col87[6];
   data_col87[8] <= data_col87[7];
   data_col87[9] <= data_col87[8];
   data_col87[10] <= data_col87[9];
   data_col87[11] <= data_col87[10];
   data_col87[12] <= data_col87[11];
   data_col87[13] <= data_col87[12];
   data_col87[14] <= data_col87[13];
   data_col87[15] <= data_col87[14];
   data_col87[16] <= data_col87[15];
   data_col87[17] <= data_col87[16];
   data_col87[18] <= data_col87[17];
   data_col87[19] <= data_col87[18];
   data_col87[20] <= data_col87[19];
   data_col87[21] <= data_col87[20];
   data_col87[22] <= data_col87[21];
   data_col87[23] <= data_col87[22];
   data_col87[24] <= data_col87[23];
   data_col87[25] <= data_col87[24];
   data_col87[26] <= data_col87[25];
   data_col87[27] <= data_col87[26];
   data_col87[28] <= data_col87[27];
   data_col87[29] <= data_col87[28];
   data_col87[30] <= data_col87[29];
   data_col87[31] <= data_col87[30];
   data_col87[32] <= data_col87[31];
   data_col87[33] <= data_col87[32];
   data_col87[34] <= data_col87[33];
   data_col87[35] <= data_col87[34];
   data_col87[36] <= data_col87[35];
   data_col87[37] <= data_col87[36];
   data_col87[38] <= data_col87[37];
   data_col87[39] <= data_col87[38];
   data_col87[40] <= data_col87[39];
   data_col87[41] <= data_col87[40];
   data_col87[42] <= data_col87[41];
   data_col87[43] <= data_col87[42];
   data_col87[44] <= data_col87[43];
   data_col87[45] <= data_col87[44];
   data_col87[46] <= data_col87[45];
   data_col87[47] <= data_col87[46];
   data_col87[48] <= data_col87[47];
   data_col87[49] <= data_col87[48];
   data_col87[50] <= data_col87[49];
   data_col87[51] <= data_col87[50];
   data_col87[52] <= data_col87[51];
   data_col87[53] <= data_col87[52];
   data_col87[54] <= data_col87[53];
   data_col87[55] <= data_col87[54];
   data_col87[56] <= data_col87[55];
   data_col87[57] <= data_col87[56];
   data_col87[58] <= data_col87[57];
   data_col87[59] <= data_col87[58];
   data_col87[60] <= data_col87[59];
   data_col87[61] <= data_col87[60];
   data_col87[62] <= data_col87[61];
   data_col87[63] <= data_col87[62];
   data_col87[64] <= data_col87[63];
   data_col87[65] <= data_col87[64];
   data_col87[66] <= data_col87[65];
   data_col87[67] <= data_col87[66];
   data_col87[68] <= data_col87[67];
   data_col87[69] <= data_col87[68];
   data_col87[70] <= data_col87[69];
   data_col87[71] <= data_col87[70];
   data_col87[72] <= data_col87[71];
   data_col87[73] <= data_col87[72];
   data_col87[74] <= data_col87[73];
   data_col87[75] <= data_col87[74];
   data_col87[76] <= data_col87[75];
   data_col87[77] <= data_col87[76];
   data_col87[78] <= data_col87[77];
   data_col87[79] <= data_col87[78];
   data_col87[80] <= data_col87[79];
   data_col87[81] <= data_col87[80];
   data_col87[82] <= data_col87[81];
   data_col87[83] <= data_col87[82];
   data_col87[84] <= data_col87[83];
   data_col87[85] <= data_col87[84];
   data_col87[86] <= data_col87[85];
   data_col87[87] <= data_col87[86];

   data_col88[1] <= data[77];
   data_col88[2] <= data_col88[1];
   data_col88[3] <= data_col88[2];
   data_col88[4] <= data_col88[3];
   data_col88[5] <= data_col88[4];
   data_col88[6] <= data_col88[5];
   data_col88[7] <= data_col88[6];
   data_col88[8] <= data_col88[7];
   data_col88[9] <= data_col88[8];
   data_col88[10] <= data_col88[9];
   data_col88[11] <= data_col88[10];
   data_col88[12] <= data_col88[11];
   data_col88[13] <= data_col88[12];
   data_col88[14] <= data_col88[13];
   data_col88[15] <= data_col88[14];
   data_col88[16] <= data_col88[15];
   data_col88[17] <= data_col88[16];
   data_col88[18] <= data_col88[17];
   data_col88[19] <= data_col88[18];
   data_col88[20] <= data_col88[19];
   data_col88[21] <= data_col88[20];
   data_col88[22] <= data_col88[21];
   data_col88[23] <= data_col88[22];
   data_col88[24] <= data_col88[23];
   data_col88[25] <= data_col88[24];
   data_col88[26] <= data_col88[25];
   data_col88[27] <= data_col88[26];
   data_col88[28] <= data_col88[27];
   data_col88[29] <= data_col88[28];
   data_col88[30] <= data_col88[29];
   data_col88[31] <= data_col88[30];
   data_col88[32] <= data_col88[31];
   data_col88[33] <= data_col88[32];
   data_col88[34] <= data_col88[33];
   data_col88[35] <= data_col88[34];
   data_col88[36] <= data_col88[35];
   data_col88[37] <= data_col88[36];
   data_col88[38] <= data_col88[37];
   data_col88[39] <= data_col88[38];
   data_col88[40] <= data_col88[39];
   data_col88[41] <= data_col88[40];
   data_col88[42] <= data_col88[41];
   data_col88[43] <= data_col88[42];
   data_col88[44] <= data_col88[43];
   data_col88[45] <= data_col88[44];
   data_col88[46] <= data_col88[45];
   data_col88[47] <= data_col88[46];
   data_col88[48] <= data_col88[47];
   data_col88[49] <= data_col88[48];
   data_col88[50] <= data_col88[49];
   data_col88[51] <= data_col88[50];
   data_col88[52] <= data_col88[51];
   data_col88[53] <= data_col88[52];
   data_col88[54] <= data_col88[53];
   data_col88[55] <= data_col88[54];
   data_col88[56] <= data_col88[55];
   data_col88[57] <= data_col88[56];
   data_col88[58] <= data_col88[57];
   data_col88[59] <= data_col88[58];
   data_col88[60] <= data_col88[59];
   data_col88[61] <= data_col88[60];
   data_col88[62] <= data_col88[61];
   data_col88[63] <= data_col88[62];
   data_col88[64] <= data_col88[63];
   data_col88[65] <= data_col88[64];
   data_col88[66] <= data_col88[65];
   data_col88[67] <= data_col88[66];
   data_col88[68] <= data_col88[67];
   data_col88[69] <= data_col88[68];
   data_col88[70] <= data_col88[69];
   data_col88[71] <= data_col88[70];
   data_col88[72] <= data_col88[71];
   data_col88[73] <= data_col88[72];
   data_col88[74] <= data_col88[73];
   data_col88[75] <= data_col88[74];
   data_col88[76] <= data_col88[75];
   data_col88[77] <= data_col88[76];
   data_col88[78] <= data_col88[77];
   data_col88[79] <= data_col88[78];
   data_col88[80] <= data_col88[79];
   data_col88[81] <= data_col88[80];
   data_col88[82] <= data_col88[81];
   data_col88[83] <= data_col88[82];
   data_col88[84] <= data_col88[83];
   data_col88[85] <= data_col88[84];
   data_col88[86] <= data_col88[85];
   data_col88[87] <= data_col88[86];
   data_col88[88] <= data_col88[87];

   data_col89[1] <= data[76];
   data_col89[2] <= data_col89[1];
   data_col89[3] <= data_col89[2];
   data_col89[4] <= data_col89[3];
   data_col89[5] <= data_col89[4];
   data_col89[6] <= data_col89[5];
   data_col89[7] <= data_col89[6];
   data_col89[8] <= data_col89[7];
   data_col89[9] <= data_col89[8];
   data_col89[10] <= data_col89[9];
   data_col89[11] <= data_col89[10];
   data_col89[12] <= data_col89[11];
   data_col89[13] <= data_col89[12];
   data_col89[14] <= data_col89[13];
   data_col89[15] <= data_col89[14];
   data_col89[16] <= data_col89[15];
   data_col89[17] <= data_col89[16];
   data_col89[18] <= data_col89[17];
   data_col89[19] <= data_col89[18];
   data_col89[20] <= data_col89[19];
   data_col89[21] <= data_col89[20];
   data_col89[22] <= data_col89[21];
   data_col89[23] <= data_col89[22];
   data_col89[24] <= data_col89[23];
   data_col89[25] <= data_col89[24];
   data_col89[26] <= data_col89[25];
   data_col89[27] <= data_col89[26];
   data_col89[28] <= data_col89[27];
   data_col89[29] <= data_col89[28];
   data_col89[30] <= data_col89[29];
   data_col89[31] <= data_col89[30];
   data_col89[32] <= data_col89[31];
   data_col89[33] <= data_col89[32];
   data_col89[34] <= data_col89[33];
   data_col89[35] <= data_col89[34];
   data_col89[36] <= data_col89[35];
   data_col89[37] <= data_col89[36];
   data_col89[38] <= data_col89[37];
   data_col89[39] <= data_col89[38];
   data_col89[40] <= data_col89[39];
   data_col89[41] <= data_col89[40];
   data_col89[42] <= data_col89[41];
   data_col89[43] <= data_col89[42];
   data_col89[44] <= data_col89[43];
   data_col89[45] <= data_col89[44];
   data_col89[46] <= data_col89[45];
   data_col89[47] <= data_col89[46];
   data_col89[48] <= data_col89[47];
   data_col89[49] <= data_col89[48];
   data_col89[50] <= data_col89[49];
   data_col89[51] <= data_col89[50];
   data_col89[52] <= data_col89[51];
   data_col89[53] <= data_col89[52];
   data_col89[54] <= data_col89[53];
   data_col89[55] <= data_col89[54];
   data_col89[56] <= data_col89[55];
   data_col89[57] <= data_col89[56];
   data_col89[58] <= data_col89[57];
   data_col89[59] <= data_col89[58];
   data_col89[60] <= data_col89[59];
   data_col89[61] <= data_col89[60];
   data_col89[62] <= data_col89[61];
   data_col89[63] <= data_col89[62];
   data_col89[64] <= data_col89[63];
   data_col89[65] <= data_col89[64];
   data_col89[66] <= data_col89[65];
   data_col89[67] <= data_col89[66];
   data_col89[68] <= data_col89[67];
   data_col89[69] <= data_col89[68];
   data_col89[70] <= data_col89[69];
   data_col89[71] <= data_col89[70];
   data_col89[72] <= data_col89[71];
   data_col89[73] <= data_col89[72];
   data_col89[74] <= data_col89[73];
   data_col89[75] <= data_col89[74];
   data_col89[76] <= data_col89[75];
   data_col89[77] <= data_col89[76];
   data_col89[78] <= data_col89[77];
   data_col89[79] <= data_col89[78];
   data_col89[80] <= data_col89[79];
   data_col89[81] <= data_col89[80];
   data_col89[82] <= data_col89[81];
   data_col89[83] <= data_col89[82];
   data_col89[84] <= data_col89[83];
   data_col89[85] <= data_col89[84];
   data_col89[86] <= data_col89[85];
   data_col89[87] <= data_col89[86];
   data_col89[88] <= data_col89[87];
   data_col89[89] <= data_col89[88];

   data_col90[1] <= data[75];
   data_col90[2] <= data_col90[1];
   data_col90[3] <= data_col90[2];
   data_col90[4] <= data_col90[3];
   data_col90[5] <= data_col90[4];
   data_col90[6] <= data_col90[5];
   data_col90[7] <= data_col90[6];
   data_col90[8] <= data_col90[7];
   data_col90[9] <= data_col90[8];
   data_col90[10] <= data_col90[9];
   data_col90[11] <= data_col90[10];
   data_col90[12] <= data_col90[11];
   data_col90[13] <= data_col90[12];
   data_col90[14] <= data_col90[13];
   data_col90[15] <= data_col90[14];
   data_col90[16] <= data_col90[15];
   data_col90[17] <= data_col90[16];
   data_col90[18] <= data_col90[17];
   data_col90[19] <= data_col90[18];
   data_col90[20] <= data_col90[19];
   data_col90[21] <= data_col90[20];
   data_col90[22] <= data_col90[21];
   data_col90[23] <= data_col90[22];
   data_col90[24] <= data_col90[23];
   data_col90[25] <= data_col90[24];
   data_col90[26] <= data_col90[25];
   data_col90[27] <= data_col90[26];
   data_col90[28] <= data_col90[27];
   data_col90[29] <= data_col90[28];
   data_col90[30] <= data_col90[29];
   data_col90[31] <= data_col90[30];
   data_col90[32] <= data_col90[31];
   data_col90[33] <= data_col90[32];
   data_col90[34] <= data_col90[33];
   data_col90[35] <= data_col90[34];
   data_col90[36] <= data_col90[35];
   data_col90[37] <= data_col90[36];
   data_col90[38] <= data_col90[37];
   data_col90[39] <= data_col90[38];
   data_col90[40] <= data_col90[39];
   data_col90[41] <= data_col90[40];
   data_col90[42] <= data_col90[41];
   data_col90[43] <= data_col90[42];
   data_col90[44] <= data_col90[43];
   data_col90[45] <= data_col90[44];
   data_col90[46] <= data_col90[45];
   data_col90[47] <= data_col90[46];
   data_col90[48] <= data_col90[47];
   data_col90[49] <= data_col90[48];
   data_col90[50] <= data_col90[49];
   data_col90[51] <= data_col90[50];
   data_col90[52] <= data_col90[51];
   data_col90[53] <= data_col90[52];
   data_col90[54] <= data_col90[53];
   data_col90[55] <= data_col90[54];
   data_col90[56] <= data_col90[55];
   data_col90[57] <= data_col90[56];
   data_col90[58] <= data_col90[57];
   data_col90[59] <= data_col90[58];
   data_col90[60] <= data_col90[59];
   data_col90[61] <= data_col90[60];
   data_col90[62] <= data_col90[61];
   data_col90[63] <= data_col90[62];
   data_col90[64] <= data_col90[63];
   data_col90[65] <= data_col90[64];
   data_col90[66] <= data_col90[65];
   data_col90[67] <= data_col90[66];
   data_col90[68] <= data_col90[67];
   data_col90[69] <= data_col90[68];
   data_col90[70] <= data_col90[69];
   data_col90[71] <= data_col90[70];
   data_col90[72] <= data_col90[71];
   data_col90[73] <= data_col90[72];
   data_col90[74] <= data_col90[73];
   data_col90[75] <= data_col90[74];
   data_col90[76] <= data_col90[75];
   data_col90[77] <= data_col90[76];
   data_col90[78] <= data_col90[77];
   data_col90[79] <= data_col90[78];
   data_col90[80] <= data_col90[79];
   data_col90[81] <= data_col90[80];
   data_col90[82] <= data_col90[81];
   data_col90[83] <= data_col90[82];
   data_col90[84] <= data_col90[83];
   data_col90[85] <= data_col90[84];
   data_col90[86] <= data_col90[85];
   data_col90[87] <= data_col90[86];
   data_col90[88] <= data_col90[87];
   data_col90[89] <= data_col90[88];
   data_col90[90] <= data_col90[89];

   data_col91[1] <= data[74];
   data_col91[2] <= data_col91[1];
   data_col91[3] <= data_col91[2];
   data_col91[4] <= data_col91[3];
   data_col91[5] <= data_col91[4];
   data_col91[6] <= data_col91[5];
   data_col91[7] <= data_col91[6];
   data_col91[8] <= data_col91[7];
   data_col91[9] <= data_col91[8];
   data_col91[10] <= data_col91[9];
   data_col91[11] <= data_col91[10];
   data_col91[12] <= data_col91[11];
   data_col91[13] <= data_col91[12];
   data_col91[14] <= data_col91[13];
   data_col91[15] <= data_col91[14];
   data_col91[16] <= data_col91[15];
   data_col91[17] <= data_col91[16];
   data_col91[18] <= data_col91[17];
   data_col91[19] <= data_col91[18];
   data_col91[20] <= data_col91[19];
   data_col91[21] <= data_col91[20];
   data_col91[22] <= data_col91[21];
   data_col91[23] <= data_col91[22];
   data_col91[24] <= data_col91[23];
   data_col91[25] <= data_col91[24];
   data_col91[26] <= data_col91[25];
   data_col91[27] <= data_col91[26];
   data_col91[28] <= data_col91[27];
   data_col91[29] <= data_col91[28];
   data_col91[30] <= data_col91[29];
   data_col91[31] <= data_col91[30];
   data_col91[32] <= data_col91[31];
   data_col91[33] <= data_col91[32];
   data_col91[34] <= data_col91[33];
   data_col91[35] <= data_col91[34];
   data_col91[36] <= data_col91[35];
   data_col91[37] <= data_col91[36];
   data_col91[38] <= data_col91[37];
   data_col91[39] <= data_col91[38];
   data_col91[40] <= data_col91[39];
   data_col91[41] <= data_col91[40];
   data_col91[42] <= data_col91[41];
   data_col91[43] <= data_col91[42];
   data_col91[44] <= data_col91[43];
   data_col91[45] <= data_col91[44];
   data_col91[46] <= data_col91[45];
   data_col91[47] <= data_col91[46];
   data_col91[48] <= data_col91[47];
   data_col91[49] <= data_col91[48];
   data_col91[50] <= data_col91[49];
   data_col91[51] <= data_col91[50];
   data_col91[52] <= data_col91[51];
   data_col91[53] <= data_col91[52];
   data_col91[54] <= data_col91[53];
   data_col91[55] <= data_col91[54];
   data_col91[56] <= data_col91[55];
   data_col91[57] <= data_col91[56];
   data_col91[58] <= data_col91[57];
   data_col91[59] <= data_col91[58];
   data_col91[60] <= data_col91[59];
   data_col91[61] <= data_col91[60];
   data_col91[62] <= data_col91[61];
   data_col91[63] <= data_col91[62];
   data_col91[64] <= data_col91[63];
   data_col91[65] <= data_col91[64];
   data_col91[66] <= data_col91[65];
   data_col91[67] <= data_col91[66];
   data_col91[68] <= data_col91[67];
   data_col91[69] <= data_col91[68];
   data_col91[70] <= data_col91[69];
   data_col91[71] <= data_col91[70];
   data_col91[72] <= data_col91[71];
   data_col91[73] <= data_col91[72];
   data_col91[74] <= data_col91[73];
   data_col91[75] <= data_col91[74];
   data_col91[76] <= data_col91[75];
   data_col91[77] <= data_col91[76];
   data_col91[78] <= data_col91[77];
   data_col91[79] <= data_col91[78];
   data_col91[80] <= data_col91[79];
   data_col91[81] <= data_col91[80];
   data_col91[82] <= data_col91[81];
   data_col91[83] <= data_col91[82];
   data_col91[84] <= data_col91[83];
   data_col91[85] <= data_col91[84];
   data_col91[86] <= data_col91[85];
   data_col91[87] <= data_col91[86];
   data_col91[88] <= data_col91[87];
   data_col91[89] <= data_col91[88];
   data_col91[90] <= data_col91[89];
   data_col91[91] <= data_col91[90];

   data_col92[1] <= data[73];
   data_col92[2] <= data_col92[1];
   data_col92[3] <= data_col92[2];
   data_col92[4] <= data_col92[3];
   data_col92[5] <= data_col92[4];
   data_col92[6] <= data_col92[5];
   data_col92[7] <= data_col92[6];
   data_col92[8] <= data_col92[7];
   data_col92[9] <= data_col92[8];
   data_col92[10] <= data_col92[9];
   data_col92[11] <= data_col92[10];
   data_col92[12] <= data_col92[11];
   data_col92[13] <= data_col92[12];
   data_col92[14] <= data_col92[13];
   data_col92[15] <= data_col92[14];
   data_col92[16] <= data_col92[15];
   data_col92[17] <= data_col92[16];
   data_col92[18] <= data_col92[17];
   data_col92[19] <= data_col92[18];
   data_col92[20] <= data_col92[19];
   data_col92[21] <= data_col92[20];
   data_col92[22] <= data_col92[21];
   data_col92[23] <= data_col92[22];
   data_col92[24] <= data_col92[23];
   data_col92[25] <= data_col92[24];
   data_col92[26] <= data_col92[25];
   data_col92[27] <= data_col92[26];
   data_col92[28] <= data_col92[27];
   data_col92[29] <= data_col92[28];
   data_col92[30] <= data_col92[29];
   data_col92[31] <= data_col92[30];
   data_col92[32] <= data_col92[31];
   data_col92[33] <= data_col92[32];
   data_col92[34] <= data_col92[33];
   data_col92[35] <= data_col92[34];
   data_col92[36] <= data_col92[35];
   data_col92[37] <= data_col92[36];
   data_col92[38] <= data_col92[37];
   data_col92[39] <= data_col92[38];
   data_col92[40] <= data_col92[39];
   data_col92[41] <= data_col92[40];
   data_col92[42] <= data_col92[41];
   data_col92[43] <= data_col92[42];
   data_col92[44] <= data_col92[43];
   data_col92[45] <= data_col92[44];
   data_col92[46] <= data_col92[45];
   data_col92[47] <= data_col92[46];
   data_col92[48] <= data_col92[47];
   data_col92[49] <= data_col92[48];
   data_col92[50] <= data_col92[49];
   data_col92[51] <= data_col92[50];
   data_col92[52] <= data_col92[51];
   data_col92[53] <= data_col92[52];
   data_col92[54] <= data_col92[53];
   data_col92[55] <= data_col92[54];
   data_col92[56] <= data_col92[55];
   data_col92[57] <= data_col92[56];
   data_col92[58] <= data_col92[57];
   data_col92[59] <= data_col92[58];
   data_col92[60] <= data_col92[59];
   data_col92[61] <= data_col92[60];
   data_col92[62] <= data_col92[61];
   data_col92[63] <= data_col92[62];
   data_col92[64] <= data_col92[63];
   data_col92[65] <= data_col92[64];
   data_col92[66] <= data_col92[65];
   data_col92[67] <= data_col92[66];
   data_col92[68] <= data_col92[67];
   data_col92[69] <= data_col92[68];
   data_col92[70] <= data_col92[69];
   data_col92[71] <= data_col92[70];
   data_col92[72] <= data_col92[71];
   data_col92[73] <= data_col92[72];
   data_col92[74] <= data_col92[73];
   data_col92[75] <= data_col92[74];
   data_col92[76] <= data_col92[75];
   data_col92[77] <= data_col92[76];
   data_col92[78] <= data_col92[77];
   data_col92[79] <= data_col92[78];
   data_col92[80] <= data_col92[79];
   data_col92[81] <= data_col92[80];
   data_col92[82] <= data_col92[81];
   data_col92[83] <= data_col92[82];
   data_col92[84] <= data_col92[83];
   data_col92[85] <= data_col92[84];
   data_col92[86] <= data_col92[85];
   data_col92[87] <= data_col92[86];
   data_col92[88] <= data_col92[87];
   data_col92[89] <= data_col92[88];
   data_col92[90] <= data_col92[89];
   data_col92[91] <= data_col92[90];
   data_col92[92] <= data_col92[91];

   data_col93[1] <= data[72];
   data_col93[2] <= data_col93[1];
   data_col93[3] <= data_col93[2];
   data_col93[4] <= data_col93[3];
   data_col93[5] <= data_col93[4];
   data_col93[6] <= data_col93[5];
   data_col93[7] <= data_col93[6];
   data_col93[8] <= data_col93[7];
   data_col93[9] <= data_col93[8];
   data_col93[10] <= data_col93[9];
   data_col93[11] <= data_col93[10];
   data_col93[12] <= data_col93[11];
   data_col93[13] <= data_col93[12];
   data_col93[14] <= data_col93[13];
   data_col93[15] <= data_col93[14];
   data_col93[16] <= data_col93[15];
   data_col93[17] <= data_col93[16];
   data_col93[18] <= data_col93[17];
   data_col93[19] <= data_col93[18];
   data_col93[20] <= data_col93[19];
   data_col93[21] <= data_col93[20];
   data_col93[22] <= data_col93[21];
   data_col93[23] <= data_col93[22];
   data_col93[24] <= data_col93[23];
   data_col93[25] <= data_col93[24];
   data_col93[26] <= data_col93[25];
   data_col93[27] <= data_col93[26];
   data_col93[28] <= data_col93[27];
   data_col93[29] <= data_col93[28];
   data_col93[30] <= data_col93[29];
   data_col93[31] <= data_col93[30];
   data_col93[32] <= data_col93[31];
   data_col93[33] <= data_col93[32];
   data_col93[34] <= data_col93[33];
   data_col93[35] <= data_col93[34];
   data_col93[36] <= data_col93[35];
   data_col93[37] <= data_col93[36];
   data_col93[38] <= data_col93[37];
   data_col93[39] <= data_col93[38];
   data_col93[40] <= data_col93[39];
   data_col93[41] <= data_col93[40];
   data_col93[42] <= data_col93[41];
   data_col93[43] <= data_col93[42];
   data_col93[44] <= data_col93[43];
   data_col93[45] <= data_col93[44];
   data_col93[46] <= data_col93[45];
   data_col93[47] <= data_col93[46];
   data_col93[48] <= data_col93[47];
   data_col93[49] <= data_col93[48];
   data_col93[50] <= data_col93[49];
   data_col93[51] <= data_col93[50];
   data_col93[52] <= data_col93[51];
   data_col93[53] <= data_col93[52];
   data_col93[54] <= data_col93[53];
   data_col93[55] <= data_col93[54];
   data_col93[56] <= data_col93[55];
   data_col93[57] <= data_col93[56];
   data_col93[58] <= data_col93[57];
   data_col93[59] <= data_col93[58];
   data_col93[60] <= data_col93[59];
   data_col93[61] <= data_col93[60];
   data_col93[62] <= data_col93[61];
   data_col93[63] <= data_col93[62];
   data_col93[64] <= data_col93[63];
   data_col93[65] <= data_col93[64];
   data_col93[66] <= data_col93[65];
   data_col93[67] <= data_col93[66];
   data_col93[68] <= data_col93[67];
   data_col93[69] <= data_col93[68];
   data_col93[70] <= data_col93[69];
   data_col93[71] <= data_col93[70];
   data_col93[72] <= data_col93[71];
   data_col93[73] <= data_col93[72];
   data_col93[74] <= data_col93[73];
   data_col93[75] <= data_col93[74];
   data_col93[76] <= data_col93[75];
   data_col93[77] <= data_col93[76];
   data_col93[78] <= data_col93[77];
   data_col93[79] <= data_col93[78];
   data_col93[80] <= data_col93[79];
   data_col93[81] <= data_col93[80];
   data_col93[82] <= data_col93[81];
   data_col93[83] <= data_col93[82];
   data_col93[84] <= data_col93[83];
   data_col93[85] <= data_col93[84];
   data_col93[86] <= data_col93[85];
   data_col93[87] <= data_col93[86];
   data_col93[88] <= data_col93[87];
   data_col93[89] <= data_col93[88];
   data_col93[90] <= data_col93[89];
   data_col93[91] <= data_col93[90];
   data_col93[92] <= data_col93[91];
   data_col93[93] <= data_col93[92];

   data_col94[1] <= data[71];
   data_col94[2] <= data_col94[1];
   data_col94[3] <= data_col94[2];
   data_col94[4] <= data_col94[3];
   data_col94[5] <= data_col94[4];
   data_col94[6] <= data_col94[5];
   data_col94[7] <= data_col94[6];
   data_col94[8] <= data_col94[7];
   data_col94[9] <= data_col94[8];
   data_col94[10] <= data_col94[9];
   data_col94[11] <= data_col94[10];
   data_col94[12] <= data_col94[11];
   data_col94[13] <= data_col94[12];
   data_col94[14] <= data_col94[13];
   data_col94[15] <= data_col94[14];
   data_col94[16] <= data_col94[15];
   data_col94[17] <= data_col94[16];
   data_col94[18] <= data_col94[17];
   data_col94[19] <= data_col94[18];
   data_col94[20] <= data_col94[19];
   data_col94[21] <= data_col94[20];
   data_col94[22] <= data_col94[21];
   data_col94[23] <= data_col94[22];
   data_col94[24] <= data_col94[23];
   data_col94[25] <= data_col94[24];
   data_col94[26] <= data_col94[25];
   data_col94[27] <= data_col94[26];
   data_col94[28] <= data_col94[27];
   data_col94[29] <= data_col94[28];
   data_col94[30] <= data_col94[29];
   data_col94[31] <= data_col94[30];
   data_col94[32] <= data_col94[31];
   data_col94[33] <= data_col94[32];
   data_col94[34] <= data_col94[33];
   data_col94[35] <= data_col94[34];
   data_col94[36] <= data_col94[35];
   data_col94[37] <= data_col94[36];
   data_col94[38] <= data_col94[37];
   data_col94[39] <= data_col94[38];
   data_col94[40] <= data_col94[39];
   data_col94[41] <= data_col94[40];
   data_col94[42] <= data_col94[41];
   data_col94[43] <= data_col94[42];
   data_col94[44] <= data_col94[43];
   data_col94[45] <= data_col94[44];
   data_col94[46] <= data_col94[45];
   data_col94[47] <= data_col94[46];
   data_col94[48] <= data_col94[47];
   data_col94[49] <= data_col94[48];
   data_col94[50] <= data_col94[49];
   data_col94[51] <= data_col94[50];
   data_col94[52] <= data_col94[51];
   data_col94[53] <= data_col94[52];
   data_col94[54] <= data_col94[53];
   data_col94[55] <= data_col94[54];
   data_col94[56] <= data_col94[55];
   data_col94[57] <= data_col94[56];
   data_col94[58] <= data_col94[57];
   data_col94[59] <= data_col94[58];
   data_col94[60] <= data_col94[59];
   data_col94[61] <= data_col94[60];
   data_col94[62] <= data_col94[61];
   data_col94[63] <= data_col94[62];
   data_col94[64] <= data_col94[63];
   data_col94[65] <= data_col94[64];
   data_col94[66] <= data_col94[65];
   data_col94[67] <= data_col94[66];
   data_col94[68] <= data_col94[67];
   data_col94[69] <= data_col94[68];
   data_col94[70] <= data_col94[69];
   data_col94[71] <= data_col94[70];
   data_col94[72] <= data_col94[71];
   data_col94[73] <= data_col94[72];
   data_col94[74] <= data_col94[73];
   data_col94[75] <= data_col94[74];
   data_col94[76] <= data_col94[75];
   data_col94[77] <= data_col94[76];
   data_col94[78] <= data_col94[77];
   data_col94[79] <= data_col94[78];
   data_col94[80] <= data_col94[79];
   data_col94[81] <= data_col94[80];
   data_col94[82] <= data_col94[81];
   data_col94[83] <= data_col94[82];
   data_col94[84] <= data_col94[83];
   data_col94[85] <= data_col94[84];
   data_col94[86] <= data_col94[85];
   data_col94[87] <= data_col94[86];
   data_col94[88] <= data_col94[87];
   data_col94[89] <= data_col94[88];
   data_col94[90] <= data_col94[89];
   data_col94[91] <= data_col94[90];
   data_col94[92] <= data_col94[91];
   data_col94[93] <= data_col94[92];
   data_col94[94] <= data_col94[93];

   data_col95[1] <= data[70];
   data_col95[2] <= data_col95[1];
   data_col95[3] <= data_col95[2];
   data_col95[4] <= data_col95[3];
   data_col95[5] <= data_col95[4];
   data_col95[6] <= data_col95[5];
   data_col95[7] <= data_col95[6];
   data_col95[8] <= data_col95[7];
   data_col95[9] <= data_col95[8];
   data_col95[10] <= data_col95[9];
   data_col95[11] <= data_col95[10];
   data_col95[12] <= data_col95[11];
   data_col95[13] <= data_col95[12];
   data_col95[14] <= data_col95[13];
   data_col95[15] <= data_col95[14];
   data_col95[16] <= data_col95[15];
   data_col95[17] <= data_col95[16];
   data_col95[18] <= data_col95[17];
   data_col95[19] <= data_col95[18];
   data_col95[20] <= data_col95[19];
   data_col95[21] <= data_col95[20];
   data_col95[22] <= data_col95[21];
   data_col95[23] <= data_col95[22];
   data_col95[24] <= data_col95[23];
   data_col95[25] <= data_col95[24];
   data_col95[26] <= data_col95[25];
   data_col95[27] <= data_col95[26];
   data_col95[28] <= data_col95[27];
   data_col95[29] <= data_col95[28];
   data_col95[30] <= data_col95[29];
   data_col95[31] <= data_col95[30];
   data_col95[32] <= data_col95[31];
   data_col95[33] <= data_col95[32];
   data_col95[34] <= data_col95[33];
   data_col95[35] <= data_col95[34];
   data_col95[36] <= data_col95[35];
   data_col95[37] <= data_col95[36];
   data_col95[38] <= data_col95[37];
   data_col95[39] <= data_col95[38];
   data_col95[40] <= data_col95[39];
   data_col95[41] <= data_col95[40];
   data_col95[42] <= data_col95[41];
   data_col95[43] <= data_col95[42];
   data_col95[44] <= data_col95[43];
   data_col95[45] <= data_col95[44];
   data_col95[46] <= data_col95[45];
   data_col95[47] <= data_col95[46];
   data_col95[48] <= data_col95[47];
   data_col95[49] <= data_col95[48];
   data_col95[50] <= data_col95[49];
   data_col95[51] <= data_col95[50];
   data_col95[52] <= data_col95[51];
   data_col95[53] <= data_col95[52];
   data_col95[54] <= data_col95[53];
   data_col95[55] <= data_col95[54];
   data_col95[56] <= data_col95[55];
   data_col95[57] <= data_col95[56];
   data_col95[58] <= data_col95[57];
   data_col95[59] <= data_col95[58];
   data_col95[60] <= data_col95[59];
   data_col95[61] <= data_col95[60];
   data_col95[62] <= data_col95[61];
   data_col95[63] <= data_col95[62];
   data_col95[64] <= data_col95[63];
   data_col95[65] <= data_col95[64];
   data_col95[66] <= data_col95[65];
   data_col95[67] <= data_col95[66];
   data_col95[68] <= data_col95[67];
   data_col95[69] <= data_col95[68];
   data_col95[70] <= data_col95[69];
   data_col95[71] <= data_col95[70];
   data_col95[72] <= data_col95[71];
   data_col95[73] <= data_col95[72];
   data_col95[74] <= data_col95[73];
   data_col95[75] <= data_col95[74];
   data_col95[76] <= data_col95[75];
   data_col95[77] <= data_col95[76];
   data_col95[78] <= data_col95[77];
   data_col95[79] <= data_col95[78];
   data_col95[80] <= data_col95[79];
   data_col95[81] <= data_col95[80];
   data_col95[82] <= data_col95[81];
   data_col95[83] <= data_col95[82];
   data_col95[84] <= data_col95[83];
   data_col95[85] <= data_col95[84];
   data_col95[86] <= data_col95[85];
   data_col95[87] <= data_col95[86];
   data_col95[88] <= data_col95[87];
   data_col95[89] <= data_col95[88];
   data_col95[90] <= data_col95[89];
   data_col95[91] <= data_col95[90];
   data_col95[92] <= data_col95[91];
   data_col95[93] <= data_col95[92];
   data_col95[94] <= data_col95[93];
   data_col95[95] <= data_col95[94];

   data_col96[1] <= data[69];
   data_col96[2] <= data_col96[1];
   data_col96[3] <= data_col96[2];
   data_col96[4] <= data_col96[3];
   data_col96[5] <= data_col96[4];
   data_col96[6] <= data_col96[5];
   data_col96[7] <= data_col96[6];
   data_col96[8] <= data_col96[7];
   data_col96[9] <= data_col96[8];
   data_col96[10] <= data_col96[9];
   data_col96[11] <= data_col96[10];
   data_col96[12] <= data_col96[11];
   data_col96[13] <= data_col96[12];
   data_col96[14] <= data_col96[13];
   data_col96[15] <= data_col96[14];
   data_col96[16] <= data_col96[15];
   data_col96[17] <= data_col96[16];
   data_col96[18] <= data_col96[17];
   data_col96[19] <= data_col96[18];
   data_col96[20] <= data_col96[19];
   data_col96[21] <= data_col96[20];
   data_col96[22] <= data_col96[21];
   data_col96[23] <= data_col96[22];
   data_col96[24] <= data_col96[23];
   data_col96[25] <= data_col96[24];
   data_col96[26] <= data_col96[25];
   data_col96[27] <= data_col96[26];
   data_col96[28] <= data_col96[27];
   data_col96[29] <= data_col96[28];
   data_col96[30] <= data_col96[29];
   data_col96[31] <= data_col96[30];
   data_col96[32] <= data_col96[31];
   data_col96[33] <= data_col96[32];
   data_col96[34] <= data_col96[33];
   data_col96[35] <= data_col96[34];
   data_col96[36] <= data_col96[35];
   data_col96[37] <= data_col96[36];
   data_col96[38] <= data_col96[37];
   data_col96[39] <= data_col96[38];
   data_col96[40] <= data_col96[39];
   data_col96[41] <= data_col96[40];
   data_col96[42] <= data_col96[41];
   data_col96[43] <= data_col96[42];
   data_col96[44] <= data_col96[43];
   data_col96[45] <= data_col96[44];
   data_col96[46] <= data_col96[45];
   data_col96[47] <= data_col96[46];
   data_col96[48] <= data_col96[47];
   data_col96[49] <= data_col96[48];
   data_col96[50] <= data_col96[49];
   data_col96[51] <= data_col96[50];
   data_col96[52] <= data_col96[51];
   data_col96[53] <= data_col96[52];
   data_col96[54] <= data_col96[53];
   data_col96[55] <= data_col96[54];
   data_col96[56] <= data_col96[55];
   data_col96[57] <= data_col96[56];
   data_col96[58] <= data_col96[57];
   data_col96[59] <= data_col96[58];
   data_col96[60] <= data_col96[59];
   data_col96[61] <= data_col96[60];
   data_col96[62] <= data_col96[61];
   data_col96[63] <= data_col96[62];
   data_col96[64] <= data_col96[63];
   data_col96[65] <= data_col96[64];
   data_col96[66] <= data_col96[65];
   data_col96[67] <= data_col96[66];
   data_col96[68] <= data_col96[67];
   data_col96[69] <= data_col96[68];
   data_col96[70] <= data_col96[69];
   data_col96[71] <= data_col96[70];
   data_col96[72] <= data_col96[71];
   data_col96[73] <= data_col96[72];
   data_col96[74] <= data_col96[73];
   data_col96[75] <= data_col96[74];
   data_col96[76] <= data_col96[75];
   data_col96[77] <= data_col96[76];
   data_col96[78] <= data_col96[77];
   data_col96[79] <= data_col96[78];
   data_col96[80] <= data_col96[79];
   data_col96[81] <= data_col96[80];
   data_col96[82] <= data_col96[81];
   data_col96[83] <= data_col96[82];
   data_col96[84] <= data_col96[83];
   data_col96[85] <= data_col96[84];
   data_col96[86] <= data_col96[85];
   data_col96[87] <= data_col96[86];
   data_col96[88] <= data_col96[87];
   data_col96[89] <= data_col96[88];
   data_col96[90] <= data_col96[89];
   data_col96[91] <= data_col96[90];
   data_col96[92] <= data_col96[91];
   data_col96[93] <= data_col96[92];
   data_col96[94] <= data_col96[93];
   data_col96[95] <= data_col96[94];
   data_col96[96] <= data_col96[95];

   data_col97[1] <= data[68];
   data_col97[2] <= data_col97[1];
   data_col97[3] <= data_col97[2];
   data_col97[4] <= data_col97[3];
   data_col97[5] <= data_col97[4];
   data_col97[6] <= data_col97[5];
   data_col97[7] <= data_col97[6];
   data_col97[8] <= data_col97[7];
   data_col97[9] <= data_col97[8];
   data_col97[10] <= data_col97[9];
   data_col97[11] <= data_col97[10];
   data_col97[12] <= data_col97[11];
   data_col97[13] <= data_col97[12];
   data_col97[14] <= data_col97[13];
   data_col97[15] <= data_col97[14];
   data_col97[16] <= data_col97[15];
   data_col97[17] <= data_col97[16];
   data_col97[18] <= data_col97[17];
   data_col97[19] <= data_col97[18];
   data_col97[20] <= data_col97[19];
   data_col97[21] <= data_col97[20];
   data_col97[22] <= data_col97[21];
   data_col97[23] <= data_col97[22];
   data_col97[24] <= data_col97[23];
   data_col97[25] <= data_col97[24];
   data_col97[26] <= data_col97[25];
   data_col97[27] <= data_col97[26];
   data_col97[28] <= data_col97[27];
   data_col97[29] <= data_col97[28];
   data_col97[30] <= data_col97[29];
   data_col97[31] <= data_col97[30];
   data_col97[32] <= data_col97[31];
   data_col97[33] <= data_col97[32];
   data_col97[34] <= data_col97[33];
   data_col97[35] <= data_col97[34];
   data_col97[36] <= data_col97[35];
   data_col97[37] <= data_col97[36];
   data_col97[38] <= data_col97[37];
   data_col97[39] <= data_col97[38];
   data_col97[40] <= data_col97[39];
   data_col97[41] <= data_col97[40];
   data_col97[42] <= data_col97[41];
   data_col97[43] <= data_col97[42];
   data_col97[44] <= data_col97[43];
   data_col97[45] <= data_col97[44];
   data_col97[46] <= data_col97[45];
   data_col97[47] <= data_col97[46];
   data_col97[48] <= data_col97[47];
   data_col97[49] <= data_col97[48];
   data_col97[50] <= data_col97[49];
   data_col97[51] <= data_col97[50];
   data_col97[52] <= data_col97[51];
   data_col97[53] <= data_col97[52];
   data_col97[54] <= data_col97[53];
   data_col97[55] <= data_col97[54];
   data_col97[56] <= data_col97[55];
   data_col97[57] <= data_col97[56];
   data_col97[58] <= data_col97[57];
   data_col97[59] <= data_col97[58];
   data_col97[60] <= data_col97[59];
   data_col97[61] <= data_col97[60];
   data_col97[62] <= data_col97[61];
   data_col97[63] <= data_col97[62];
   data_col97[64] <= data_col97[63];
   data_col97[65] <= data_col97[64];
   data_col97[66] <= data_col97[65];
   data_col97[67] <= data_col97[66];
   data_col97[68] <= data_col97[67];
   data_col97[69] <= data_col97[68];
   data_col97[70] <= data_col97[69];
   data_col97[71] <= data_col97[70];
   data_col97[72] <= data_col97[71];
   data_col97[73] <= data_col97[72];
   data_col97[74] <= data_col97[73];
   data_col97[75] <= data_col97[74];
   data_col97[76] <= data_col97[75];
   data_col97[77] <= data_col97[76];
   data_col97[78] <= data_col97[77];
   data_col97[79] <= data_col97[78];
   data_col97[80] <= data_col97[79];
   data_col97[81] <= data_col97[80];
   data_col97[82] <= data_col97[81];
   data_col97[83] <= data_col97[82];
   data_col97[84] <= data_col97[83];
   data_col97[85] <= data_col97[84];
   data_col97[86] <= data_col97[85];
   data_col97[87] <= data_col97[86];
   data_col97[88] <= data_col97[87];
   data_col97[89] <= data_col97[88];
   data_col97[90] <= data_col97[89];
   data_col97[91] <= data_col97[90];
   data_col97[92] <= data_col97[91];
   data_col97[93] <= data_col97[92];
   data_col97[94] <= data_col97[93];
   data_col97[95] <= data_col97[94];
   data_col97[96] <= data_col97[95];
   data_col97[97] <= data_col97[96];

   data_col98[1] <= data[67];
   data_col98[2] <= data_col98[1];
   data_col98[3] <= data_col98[2];
   data_col98[4] <= data_col98[3];
   data_col98[5] <= data_col98[4];
   data_col98[6] <= data_col98[5];
   data_col98[7] <= data_col98[6];
   data_col98[8] <= data_col98[7];
   data_col98[9] <= data_col98[8];
   data_col98[10] <= data_col98[9];
   data_col98[11] <= data_col98[10];
   data_col98[12] <= data_col98[11];
   data_col98[13] <= data_col98[12];
   data_col98[14] <= data_col98[13];
   data_col98[15] <= data_col98[14];
   data_col98[16] <= data_col98[15];
   data_col98[17] <= data_col98[16];
   data_col98[18] <= data_col98[17];
   data_col98[19] <= data_col98[18];
   data_col98[20] <= data_col98[19];
   data_col98[21] <= data_col98[20];
   data_col98[22] <= data_col98[21];
   data_col98[23] <= data_col98[22];
   data_col98[24] <= data_col98[23];
   data_col98[25] <= data_col98[24];
   data_col98[26] <= data_col98[25];
   data_col98[27] <= data_col98[26];
   data_col98[28] <= data_col98[27];
   data_col98[29] <= data_col98[28];
   data_col98[30] <= data_col98[29];
   data_col98[31] <= data_col98[30];
   data_col98[32] <= data_col98[31];
   data_col98[33] <= data_col98[32];
   data_col98[34] <= data_col98[33];
   data_col98[35] <= data_col98[34];
   data_col98[36] <= data_col98[35];
   data_col98[37] <= data_col98[36];
   data_col98[38] <= data_col98[37];
   data_col98[39] <= data_col98[38];
   data_col98[40] <= data_col98[39];
   data_col98[41] <= data_col98[40];
   data_col98[42] <= data_col98[41];
   data_col98[43] <= data_col98[42];
   data_col98[44] <= data_col98[43];
   data_col98[45] <= data_col98[44];
   data_col98[46] <= data_col98[45];
   data_col98[47] <= data_col98[46];
   data_col98[48] <= data_col98[47];
   data_col98[49] <= data_col98[48];
   data_col98[50] <= data_col98[49];
   data_col98[51] <= data_col98[50];
   data_col98[52] <= data_col98[51];
   data_col98[53] <= data_col98[52];
   data_col98[54] <= data_col98[53];
   data_col98[55] <= data_col98[54];
   data_col98[56] <= data_col98[55];
   data_col98[57] <= data_col98[56];
   data_col98[58] <= data_col98[57];
   data_col98[59] <= data_col98[58];
   data_col98[60] <= data_col98[59];
   data_col98[61] <= data_col98[60];
   data_col98[62] <= data_col98[61];
   data_col98[63] <= data_col98[62];
   data_col98[64] <= data_col98[63];
   data_col98[65] <= data_col98[64];
   data_col98[66] <= data_col98[65];
   data_col98[67] <= data_col98[66];
   data_col98[68] <= data_col98[67];
   data_col98[69] <= data_col98[68];
   data_col98[70] <= data_col98[69];
   data_col98[71] <= data_col98[70];
   data_col98[72] <= data_col98[71];
   data_col98[73] <= data_col98[72];
   data_col98[74] <= data_col98[73];
   data_col98[75] <= data_col98[74];
   data_col98[76] <= data_col98[75];
   data_col98[77] <= data_col98[76];
   data_col98[78] <= data_col98[77];
   data_col98[79] <= data_col98[78];
   data_col98[80] <= data_col98[79];
   data_col98[81] <= data_col98[80];
   data_col98[82] <= data_col98[81];
   data_col98[83] <= data_col98[82];
   data_col98[84] <= data_col98[83];
   data_col98[85] <= data_col98[84];
   data_col98[86] <= data_col98[85];
   data_col98[87] <= data_col98[86];
   data_col98[88] <= data_col98[87];
   data_col98[89] <= data_col98[88];
   data_col98[90] <= data_col98[89];
   data_col98[91] <= data_col98[90];
   data_col98[92] <= data_col98[91];
   data_col98[93] <= data_col98[92];
   data_col98[94] <= data_col98[93];
   data_col98[95] <= data_col98[94];
   data_col98[96] <= data_col98[95];
   data_col98[97] <= data_col98[96];
   data_col98[98] <= data_col98[97];

   data_col99[1] <= data[66];
   data_col99[2] <= data_col99[1];
   data_col99[3] <= data_col99[2];
   data_col99[4] <= data_col99[3];
   data_col99[5] <= data_col99[4];
   data_col99[6] <= data_col99[5];
   data_col99[7] <= data_col99[6];
   data_col99[8] <= data_col99[7];
   data_col99[9] <= data_col99[8];
   data_col99[10] <= data_col99[9];
   data_col99[11] <= data_col99[10];
   data_col99[12] <= data_col99[11];
   data_col99[13] <= data_col99[12];
   data_col99[14] <= data_col99[13];
   data_col99[15] <= data_col99[14];
   data_col99[16] <= data_col99[15];
   data_col99[17] <= data_col99[16];
   data_col99[18] <= data_col99[17];
   data_col99[19] <= data_col99[18];
   data_col99[20] <= data_col99[19];
   data_col99[21] <= data_col99[20];
   data_col99[22] <= data_col99[21];
   data_col99[23] <= data_col99[22];
   data_col99[24] <= data_col99[23];
   data_col99[25] <= data_col99[24];
   data_col99[26] <= data_col99[25];
   data_col99[27] <= data_col99[26];
   data_col99[28] <= data_col99[27];
   data_col99[29] <= data_col99[28];
   data_col99[30] <= data_col99[29];
   data_col99[31] <= data_col99[30];
   data_col99[32] <= data_col99[31];
   data_col99[33] <= data_col99[32];
   data_col99[34] <= data_col99[33];
   data_col99[35] <= data_col99[34];
   data_col99[36] <= data_col99[35];
   data_col99[37] <= data_col99[36];
   data_col99[38] <= data_col99[37];
   data_col99[39] <= data_col99[38];
   data_col99[40] <= data_col99[39];
   data_col99[41] <= data_col99[40];
   data_col99[42] <= data_col99[41];
   data_col99[43] <= data_col99[42];
   data_col99[44] <= data_col99[43];
   data_col99[45] <= data_col99[44];
   data_col99[46] <= data_col99[45];
   data_col99[47] <= data_col99[46];
   data_col99[48] <= data_col99[47];
   data_col99[49] <= data_col99[48];
   data_col99[50] <= data_col99[49];
   data_col99[51] <= data_col99[50];
   data_col99[52] <= data_col99[51];
   data_col99[53] <= data_col99[52];
   data_col99[54] <= data_col99[53];
   data_col99[55] <= data_col99[54];
   data_col99[56] <= data_col99[55];
   data_col99[57] <= data_col99[56];
   data_col99[58] <= data_col99[57];
   data_col99[59] <= data_col99[58];
   data_col99[60] <= data_col99[59];
   data_col99[61] <= data_col99[60];
   data_col99[62] <= data_col99[61];
   data_col99[63] <= data_col99[62];
   data_col99[64] <= data_col99[63];
   data_col99[65] <= data_col99[64];
   data_col99[66] <= data_col99[65];
   data_col99[67] <= data_col99[66];
   data_col99[68] <= data_col99[67];
   data_col99[69] <= data_col99[68];
   data_col99[70] <= data_col99[69];
   data_col99[71] <= data_col99[70];
   data_col99[72] <= data_col99[71];
   data_col99[73] <= data_col99[72];
   data_col99[74] <= data_col99[73];
   data_col99[75] <= data_col99[74];
   data_col99[76] <= data_col99[75];
   data_col99[77] <= data_col99[76];
   data_col99[78] <= data_col99[77];
   data_col99[79] <= data_col99[78];
   data_col99[80] <= data_col99[79];
   data_col99[81] <= data_col99[80];
   data_col99[82] <= data_col99[81];
   data_col99[83] <= data_col99[82];
   data_col99[84] <= data_col99[83];
   data_col99[85] <= data_col99[84];
   data_col99[86] <= data_col99[85];
   data_col99[87] <= data_col99[86];
   data_col99[88] <= data_col99[87];
   data_col99[89] <= data_col99[88];
   data_col99[90] <= data_col99[89];
   data_col99[91] <= data_col99[90];
   data_col99[92] <= data_col99[91];
   data_col99[93] <= data_col99[92];
   data_col99[94] <= data_col99[93];
   data_col99[95] <= data_col99[94];
   data_col99[96] <= data_col99[95];
   data_col99[97] <= data_col99[96];
   data_col99[98] <= data_col99[97];
   data_col99[99] <= data_col99[98];

   data_col100[1] <= data[65];
   data_col100[2] <= data_col100[1];
   data_col100[3] <= data_col100[2];
   data_col100[4] <= data_col100[3];
   data_col100[5] <= data_col100[4];
   data_col100[6] <= data_col100[5];
   data_col100[7] <= data_col100[6];
   data_col100[8] <= data_col100[7];
   data_col100[9] <= data_col100[8];
   data_col100[10] <= data_col100[9];
   data_col100[11] <= data_col100[10];
   data_col100[12] <= data_col100[11];
   data_col100[13] <= data_col100[12];
   data_col100[14] <= data_col100[13];
   data_col100[15] <= data_col100[14];
   data_col100[16] <= data_col100[15];
   data_col100[17] <= data_col100[16];
   data_col100[18] <= data_col100[17];
   data_col100[19] <= data_col100[18];
   data_col100[20] <= data_col100[19];
   data_col100[21] <= data_col100[20];
   data_col100[22] <= data_col100[21];
   data_col100[23] <= data_col100[22];
   data_col100[24] <= data_col100[23];
   data_col100[25] <= data_col100[24];
   data_col100[26] <= data_col100[25];
   data_col100[27] <= data_col100[26];
   data_col100[28] <= data_col100[27];
   data_col100[29] <= data_col100[28];
   data_col100[30] <= data_col100[29];
   data_col100[31] <= data_col100[30];
   data_col100[32] <= data_col100[31];
   data_col100[33] <= data_col100[32];
   data_col100[34] <= data_col100[33];
   data_col100[35] <= data_col100[34];
   data_col100[36] <= data_col100[35];
   data_col100[37] <= data_col100[36];
   data_col100[38] <= data_col100[37];
   data_col100[39] <= data_col100[38];
   data_col100[40] <= data_col100[39];
   data_col100[41] <= data_col100[40];
   data_col100[42] <= data_col100[41];
   data_col100[43] <= data_col100[42];
   data_col100[44] <= data_col100[43];
   data_col100[45] <= data_col100[44];
   data_col100[46] <= data_col100[45];
   data_col100[47] <= data_col100[46];
   data_col100[48] <= data_col100[47];
   data_col100[49] <= data_col100[48];
   data_col100[50] <= data_col100[49];
   data_col100[51] <= data_col100[50];
   data_col100[52] <= data_col100[51];
   data_col100[53] <= data_col100[52];
   data_col100[54] <= data_col100[53];
   data_col100[55] <= data_col100[54];
   data_col100[56] <= data_col100[55];
   data_col100[57] <= data_col100[56];
   data_col100[58] <= data_col100[57];
   data_col100[59] <= data_col100[58];
   data_col100[60] <= data_col100[59];
   data_col100[61] <= data_col100[60];
   data_col100[62] <= data_col100[61];
   data_col100[63] <= data_col100[62];
   data_col100[64] <= data_col100[63];
   data_col100[65] <= data_col100[64];
   data_col100[66] <= data_col100[65];
   data_col100[67] <= data_col100[66];
   data_col100[68] <= data_col100[67];
   data_col100[69] <= data_col100[68];
   data_col100[70] <= data_col100[69];
   data_col100[71] <= data_col100[70];
   data_col100[72] <= data_col100[71];
   data_col100[73] <= data_col100[72];
   data_col100[74] <= data_col100[73];
   data_col100[75] <= data_col100[74];
   data_col100[76] <= data_col100[75];
   data_col100[77] <= data_col100[76];
   data_col100[78] <= data_col100[77];
   data_col100[79] <= data_col100[78];
   data_col100[80] <= data_col100[79];
   data_col100[81] <= data_col100[80];
   data_col100[82] <= data_col100[81];
   data_col100[83] <= data_col100[82];
   data_col100[84] <= data_col100[83];
   data_col100[85] <= data_col100[84];
   data_col100[86] <= data_col100[85];
   data_col100[87] <= data_col100[86];
   data_col100[88] <= data_col100[87];
   data_col100[89] <= data_col100[88];
   data_col100[90] <= data_col100[89];
   data_col100[91] <= data_col100[90];
   data_col100[92] <= data_col100[91];
   data_col100[93] <= data_col100[92];
   data_col100[94] <= data_col100[93];
   data_col100[95] <= data_col100[94];
   data_col100[96] <= data_col100[95];
   data_col100[97] <= data_col100[96];
   data_col100[98] <= data_col100[97];
   data_col100[99] <= data_col100[98];
   data_col100[100] <= data_col100[99];

   data_col101[1] <= data[64];
   data_col101[2] <= data_col101[1];
   data_col101[3] <= data_col101[2];
   data_col101[4] <= data_col101[3];
   data_col101[5] <= data_col101[4];
   data_col101[6] <= data_col101[5];
   data_col101[7] <= data_col101[6];
   data_col101[8] <= data_col101[7];
   data_col101[9] <= data_col101[8];
   data_col101[10] <= data_col101[9];
   data_col101[11] <= data_col101[10];
   data_col101[12] <= data_col101[11];
   data_col101[13] <= data_col101[12];
   data_col101[14] <= data_col101[13];
   data_col101[15] <= data_col101[14];
   data_col101[16] <= data_col101[15];
   data_col101[17] <= data_col101[16];
   data_col101[18] <= data_col101[17];
   data_col101[19] <= data_col101[18];
   data_col101[20] <= data_col101[19];
   data_col101[21] <= data_col101[20];
   data_col101[22] <= data_col101[21];
   data_col101[23] <= data_col101[22];
   data_col101[24] <= data_col101[23];
   data_col101[25] <= data_col101[24];
   data_col101[26] <= data_col101[25];
   data_col101[27] <= data_col101[26];
   data_col101[28] <= data_col101[27];
   data_col101[29] <= data_col101[28];
   data_col101[30] <= data_col101[29];
   data_col101[31] <= data_col101[30];
   data_col101[32] <= data_col101[31];
   data_col101[33] <= data_col101[32];
   data_col101[34] <= data_col101[33];
   data_col101[35] <= data_col101[34];
   data_col101[36] <= data_col101[35];
   data_col101[37] <= data_col101[36];
   data_col101[38] <= data_col101[37];
   data_col101[39] <= data_col101[38];
   data_col101[40] <= data_col101[39];
   data_col101[41] <= data_col101[40];
   data_col101[42] <= data_col101[41];
   data_col101[43] <= data_col101[42];
   data_col101[44] <= data_col101[43];
   data_col101[45] <= data_col101[44];
   data_col101[46] <= data_col101[45];
   data_col101[47] <= data_col101[46];
   data_col101[48] <= data_col101[47];
   data_col101[49] <= data_col101[48];
   data_col101[50] <= data_col101[49];
   data_col101[51] <= data_col101[50];
   data_col101[52] <= data_col101[51];
   data_col101[53] <= data_col101[52];
   data_col101[54] <= data_col101[53];
   data_col101[55] <= data_col101[54];
   data_col101[56] <= data_col101[55];
   data_col101[57] <= data_col101[56];
   data_col101[58] <= data_col101[57];
   data_col101[59] <= data_col101[58];
   data_col101[60] <= data_col101[59];
   data_col101[61] <= data_col101[60];
   data_col101[62] <= data_col101[61];
   data_col101[63] <= data_col101[62];
   data_col101[64] <= data_col101[63];
   data_col101[65] <= data_col101[64];
   data_col101[66] <= data_col101[65];
   data_col101[67] <= data_col101[66];
   data_col101[68] <= data_col101[67];
   data_col101[69] <= data_col101[68];
   data_col101[70] <= data_col101[69];
   data_col101[71] <= data_col101[70];
   data_col101[72] <= data_col101[71];
   data_col101[73] <= data_col101[72];
   data_col101[74] <= data_col101[73];
   data_col101[75] <= data_col101[74];
   data_col101[76] <= data_col101[75];
   data_col101[77] <= data_col101[76];
   data_col101[78] <= data_col101[77];
   data_col101[79] <= data_col101[78];
   data_col101[80] <= data_col101[79];
   data_col101[81] <= data_col101[80];
   data_col101[82] <= data_col101[81];
   data_col101[83] <= data_col101[82];
   data_col101[84] <= data_col101[83];
   data_col101[85] <= data_col101[84];
   data_col101[86] <= data_col101[85];
   data_col101[87] <= data_col101[86];
   data_col101[88] <= data_col101[87];
   data_col101[89] <= data_col101[88];
   data_col101[90] <= data_col101[89];
   data_col101[91] <= data_col101[90];
   data_col101[92] <= data_col101[91];
   data_col101[93] <= data_col101[92];
   data_col101[94] <= data_col101[93];
   data_col101[95] <= data_col101[94];
   data_col101[96] <= data_col101[95];
   data_col101[97] <= data_col101[96];
   data_col101[98] <= data_col101[97];
   data_col101[99] <= data_col101[98];
   data_col101[100] <= data_col101[99];
   data_col101[101] <= data_col101[100];

   data_col102[1] <= data[63];
   data_col102[2] <= data_col102[1];
   data_col102[3] <= data_col102[2];
   data_col102[4] <= data_col102[3];
   data_col102[5] <= data_col102[4];
   data_col102[6] <= data_col102[5];
   data_col102[7] <= data_col102[6];
   data_col102[8] <= data_col102[7];
   data_col102[9] <= data_col102[8];
   data_col102[10] <= data_col102[9];
   data_col102[11] <= data_col102[10];
   data_col102[12] <= data_col102[11];
   data_col102[13] <= data_col102[12];
   data_col102[14] <= data_col102[13];
   data_col102[15] <= data_col102[14];
   data_col102[16] <= data_col102[15];
   data_col102[17] <= data_col102[16];
   data_col102[18] <= data_col102[17];
   data_col102[19] <= data_col102[18];
   data_col102[20] <= data_col102[19];
   data_col102[21] <= data_col102[20];
   data_col102[22] <= data_col102[21];
   data_col102[23] <= data_col102[22];
   data_col102[24] <= data_col102[23];
   data_col102[25] <= data_col102[24];
   data_col102[26] <= data_col102[25];
   data_col102[27] <= data_col102[26];
   data_col102[28] <= data_col102[27];
   data_col102[29] <= data_col102[28];
   data_col102[30] <= data_col102[29];
   data_col102[31] <= data_col102[30];
   data_col102[32] <= data_col102[31];
   data_col102[33] <= data_col102[32];
   data_col102[34] <= data_col102[33];
   data_col102[35] <= data_col102[34];
   data_col102[36] <= data_col102[35];
   data_col102[37] <= data_col102[36];
   data_col102[38] <= data_col102[37];
   data_col102[39] <= data_col102[38];
   data_col102[40] <= data_col102[39];
   data_col102[41] <= data_col102[40];
   data_col102[42] <= data_col102[41];
   data_col102[43] <= data_col102[42];
   data_col102[44] <= data_col102[43];
   data_col102[45] <= data_col102[44];
   data_col102[46] <= data_col102[45];
   data_col102[47] <= data_col102[46];
   data_col102[48] <= data_col102[47];
   data_col102[49] <= data_col102[48];
   data_col102[50] <= data_col102[49];
   data_col102[51] <= data_col102[50];
   data_col102[52] <= data_col102[51];
   data_col102[53] <= data_col102[52];
   data_col102[54] <= data_col102[53];
   data_col102[55] <= data_col102[54];
   data_col102[56] <= data_col102[55];
   data_col102[57] <= data_col102[56];
   data_col102[58] <= data_col102[57];
   data_col102[59] <= data_col102[58];
   data_col102[60] <= data_col102[59];
   data_col102[61] <= data_col102[60];
   data_col102[62] <= data_col102[61];
   data_col102[63] <= data_col102[62];
   data_col102[64] <= data_col102[63];
   data_col102[65] <= data_col102[64];
   data_col102[66] <= data_col102[65];
   data_col102[67] <= data_col102[66];
   data_col102[68] <= data_col102[67];
   data_col102[69] <= data_col102[68];
   data_col102[70] <= data_col102[69];
   data_col102[71] <= data_col102[70];
   data_col102[72] <= data_col102[71];
   data_col102[73] <= data_col102[72];
   data_col102[74] <= data_col102[73];
   data_col102[75] <= data_col102[74];
   data_col102[76] <= data_col102[75];
   data_col102[77] <= data_col102[76];
   data_col102[78] <= data_col102[77];
   data_col102[79] <= data_col102[78];
   data_col102[80] <= data_col102[79];
   data_col102[81] <= data_col102[80];
   data_col102[82] <= data_col102[81];
   data_col102[83] <= data_col102[82];
   data_col102[84] <= data_col102[83];
   data_col102[85] <= data_col102[84];
   data_col102[86] <= data_col102[85];
   data_col102[87] <= data_col102[86];
   data_col102[88] <= data_col102[87];
   data_col102[89] <= data_col102[88];
   data_col102[90] <= data_col102[89];
   data_col102[91] <= data_col102[90];
   data_col102[92] <= data_col102[91];
   data_col102[93] <= data_col102[92];
   data_col102[94] <= data_col102[93];
   data_col102[95] <= data_col102[94];
   data_col102[96] <= data_col102[95];
   data_col102[97] <= data_col102[96];
   data_col102[98] <= data_col102[97];
   data_col102[99] <= data_col102[98];
   data_col102[100] <= data_col102[99];
   data_col102[101] <= data_col102[100];
   data_col102[102] <= data_col102[101];

   data_col103[1] <= data[62];
   data_col103[2] <= data_col103[1];
   data_col103[3] <= data_col103[2];
   data_col103[4] <= data_col103[3];
   data_col103[5] <= data_col103[4];
   data_col103[6] <= data_col103[5];
   data_col103[7] <= data_col103[6];
   data_col103[8] <= data_col103[7];
   data_col103[9] <= data_col103[8];
   data_col103[10] <= data_col103[9];
   data_col103[11] <= data_col103[10];
   data_col103[12] <= data_col103[11];
   data_col103[13] <= data_col103[12];
   data_col103[14] <= data_col103[13];
   data_col103[15] <= data_col103[14];
   data_col103[16] <= data_col103[15];
   data_col103[17] <= data_col103[16];
   data_col103[18] <= data_col103[17];
   data_col103[19] <= data_col103[18];
   data_col103[20] <= data_col103[19];
   data_col103[21] <= data_col103[20];
   data_col103[22] <= data_col103[21];
   data_col103[23] <= data_col103[22];
   data_col103[24] <= data_col103[23];
   data_col103[25] <= data_col103[24];
   data_col103[26] <= data_col103[25];
   data_col103[27] <= data_col103[26];
   data_col103[28] <= data_col103[27];
   data_col103[29] <= data_col103[28];
   data_col103[30] <= data_col103[29];
   data_col103[31] <= data_col103[30];
   data_col103[32] <= data_col103[31];
   data_col103[33] <= data_col103[32];
   data_col103[34] <= data_col103[33];
   data_col103[35] <= data_col103[34];
   data_col103[36] <= data_col103[35];
   data_col103[37] <= data_col103[36];
   data_col103[38] <= data_col103[37];
   data_col103[39] <= data_col103[38];
   data_col103[40] <= data_col103[39];
   data_col103[41] <= data_col103[40];
   data_col103[42] <= data_col103[41];
   data_col103[43] <= data_col103[42];
   data_col103[44] <= data_col103[43];
   data_col103[45] <= data_col103[44];
   data_col103[46] <= data_col103[45];
   data_col103[47] <= data_col103[46];
   data_col103[48] <= data_col103[47];
   data_col103[49] <= data_col103[48];
   data_col103[50] <= data_col103[49];
   data_col103[51] <= data_col103[50];
   data_col103[52] <= data_col103[51];
   data_col103[53] <= data_col103[52];
   data_col103[54] <= data_col103[53];
   data_col103[55] <= data_col103[54];
   data_col103[56] <= data_col103[55];
   data_col103[57] <= data_col103[56];
   data_col103[58] <= data_col103[57];
   data_col103[59] <= data_col103[58];
   data_col103[60] <= data_col103[59];
   data_col103[61] <= data_col103[60];
   data_col103[62] <= data_col103[61];
   data_col103[63] <= data_col103[62];
   data_col103[64] <= data_col103[63];
   data_col103[65] <= data_col103[64];
   data_col103[66] <= data_col103[65];
   data_col103[67] <= data_col103[66];
   data_col103[68] <= data_col103[67];
   data_col103[69] <= data_col103[68];
   data_col103[70] <= data_col103[69];
   data_col103[71] <= data_col103[70];
   data_col103[72] <= data_col103[71];
   data_col103[73] <= data_col103[72];
   data_col103[74] <= data_col103[73];
   data_col103[75] <= data_col103[74];
   data_col103[76] <= data_col103[75];
   data_col103[77] <= data_col103[76];
   data_col103[78] <= data_col103[77];
   data_col103[79] <= data_col103[78];
   data_col103[80] <= data_col103[79];
   data_col103[81] <= data_col103[80];
   data_col103[82] <= data_col103[81];
   data_col103[83] <= data_col103[82];
   data_col103[84] <= data_col103[83];
   data_col103[85] <= data_col103[84];
   data_col103[86] <= data_col103[85];
   data_col103[87] <= data_col103[86];
   data_col103[88] <= data_col103[87];
   data_col103[89] <= data_col103[88];
   data_col103[90] <= data_col103[89];
   data_col103[91] <= data_col103[90];
   data_col103[92] <= data_col103[91];
   data_col103[93] <= data_col103[92];
   data_col103[94] <= data_col103[93];
   data_col103[95] <= data_col103[94];
   data_col103[96] <= data_col103[95];
   data_col103[97] <= data_col103[96];
   data_col103[98] <= data_col103[97];
   data_col103[99] <= data_col103[98];
   data_col103[100] <= data_col103[99];
   data_col103[101] <= data_col103[100];
   data_col103[102] <= data_col103[101];
   data_col103[103] <= data_col103[102];

   data_col104[1] <= data[61];
   data_col104[2] <= data_col104[1];
   data_col104[3] <= data_col104[2];
   data_col104[4] <= data_col104[3];
   data_col104[5] <= data_col104[4];
   data_col104[6] <= data_col104[5];
   data_col104[7] <= data_col104[6];
   data_col104[8] <= data_col104[7];
   data_col104[9] <= data_col104[8];
   data_col104[10] <= data_col104[9];
   data_col104[11] <= data_col104[10];
   data_col104[12] <= data_col104[11];
   data_col104[13] <= data_col104[12];
   data_col104[14] <= data_col104[13];
   data_col104[15] <= data_col104[14];
   data_col104[16] <= data_col104[15];
   data_col104[17] <= data_col104[16];
   data_col104[18] <= data_col104[17];
   data_col104[19] <= data_col104[18];
   data_col104[20] <= data_col104[19];
   data_col104[21] <= data_col104[20];
   data_col104[22] <= data_col104[21];
   data_col104[23] <= data_col104[22];
   data_col104[24] <= data_col104[23];
   data_col104[25] <= data_col104[24];
   data_col104[26] <= data_col104[25];
   data_col104[27] <= data_col104[26];
   data_col104[28] <= data_col104[27];
   data_col104[29] <= data_col104[28];
   data_col104[30] <= data_col104[29];
   data_col104[31] <= data_col104[30];
   data_col104[32] <= data_col104[31];
   data_col104[33] <= data_col104[32];
   data_col104[34] <= data_col104[33];
   data_col104[35] <= data_col104[34];
   data_col104[36] <= data_col104[35];
   data_col104[37] <= data_col104[36];
   data_col104[38] <= data_col104[37];
   data_col104[39] <= data_col104[38];
   data_col104[40] <= data_col104[39];
   data_col104[41] <= data_col104[40];
   data_col104[42] <= data_col104[41];
   data_col104[43] <= data_col104[42];
   data_col104[44] <= data_col104[43];
   data_col104[45] <= data_col104[44];
   data_col104[46] <= data_col104[45];
   data_col104[47] <= data_col104[46];
   data_col104[48] <= data_col104[47];
   data_col104[49] <= data_col104[48];
   data_col104[50] <= data_col104[49];
   data_col104[51] <= data_col104[50];
   data_col104[52] <= data_col104[51];
   data_col104[53] <= data_col104[52];
   data_col104[54] <= data_col104[53];
   data_col104[55] <= data_col104[54];
   data_col104[56] <= data_col104[55];
   data_col104[57] <= data_col104[56];
   data_col104[58] <= data_col104[57];
   data_col104[59] <= data_col104[58];
   data_col104[60] <= data_col104[59];
   data_col104[61] <= data_col104[60];
   data_col104[62] <= data_col104[61];
   data_col104[63] <= data_col104[62];
   data_col104[64] <= data_col104[63];
   data_col104[65] <= data_col104[64];
   data_col104[66] <= data_col104[65];
   data_col104[67] <= data_col104[66];
   data_col104[68] <= data_col104[67];
   data_col104[69] <= data_col104[68];
   data_col104[70] <= data_col104[69];
   data_col104[71] <= data_col104[70];
   data_col104[72] <= data_col104[71];
   data_col104[73] <= data_col104[72];
   data_col104[74] <= data_col104[73];
   data_col104[75] <= data_col104[74];
   data_col104[76] <= data_col104[75];
   data_col104[77] <= data_col104[76];
   data_col104[78] <= data_col104[77];
   data_col104[79] <= data_col104[78];
   data_col104[80] <= data_col104[79];
   data_col104[81] <= data_col104[80];
   data_col104[82] <= data_col104[81];
   data_col104[83] <= data_col104[82];
   data_col104[84] <= data_col104[83];
   data_col104[85] <= data_col104[84];
   data_col104[86] <= data_col104[85];
   data_col104[87] <= data_col104[86];
   data_col104[88] <= data_col104[87];
   data_col104[89] <= data_col104[88];
   data_col104[90] <= data_col104[89];
   data_col104[91] <= data_col104[90];
   data_col104[92] <= data_col104[91];
   data_col104[93] <= data_col104[92];
   data_col104[94] <= data_col104[93];
   data_col104[95] <= data_col104[94];
   data_col104[96] <= data_col104[95];
   data_col104[97] <= data_col104[96];
   data_col104[98] <= data_col104[97];
   data_col104[99] <= data_col104[98];
   data_col104[100] <= data_col104[99];
   data_col104[101] <= data_col104[100];
   data_col104[102] <= data_col104[101];
   data_col104[103] <= data_col104[102];
   data_col104[104] <= data_col104[103];

   data_col105[1] <= data[60];
   data_col105[2] <= data_col105[1];
   data_col105[3] <= data_col105[2];
   data_col105[4] <= data_col105[3];
   data_col105[5] <= data_col105[4];
   data_col105[6] <= data_col105[5];
   data_col105[7] <= data_col105[6];
   data_col105[8] <= data_col105[7];
   data_col105[9] <= data_col105[8];
   data_col105[10] <= data_col105[9];
   data_col105[11] <= data_col105[10];
   data_col105[12] <= data_col105[11];
   data_col105[13] <= data_col105[12];
   data_col105[14] <= data_col105[13];
   data_col105[15] <= data_col105[14];
   data_col105[16] <= data_col105[15];
   data_col105[17] <= data_col105[16];
   data_col105[18] <= data_col105[17];
   data_col105[19] <= data_col105[18];
   data_col105[20] <= data_col105[19];
   data_col105[21] <= data_col105[20];
   data_col105[22] <= data_col105[21];
   data_col105[23] <= data_col105[22];
   data_col105[24] <= data_col105[23];
   data_col105[25] <= data_col105[24];
   data_col105[26] <= data_col105[25];
   data_col105[27] <= data_col105[26];
   data_col105[28] <= data_col105[27];
   data_col105[29] <= data_col105[28];
   data_col105[30] <= data_col105[29];
   data_col105[31] <= data_col105[30];
   data_col105[32] <= data_col105[31];
   data_col105[33] <= data_col105[32];
   data_col105[34] <= data_col105[33];
   data_col105[35] <= data_col105[34];
   data_col105[36] <= data_col105[35];
   data_col105[37] <= data_col105[36];
   data_col105[38] <= data_col105[37];
   data_col105[39] <= data_col105[38];
   data_col105[40] <= data_col105[39];
   data_col105[41] <= data_col105[40];
   data_col105[42] <= data_col105[41];
   data_col105[43] <= data_col105[42];
   data_col105[44] <= data_col105[43];
   data_col105[45] <= data_col105[44];
   data_col105[46] <= data_col105[45];
   data_col105[47] <= data_col105[46];
   data_col105[48] <= data_col105[47];
   data_col105[49] <= data_col105[48];
   data_col105[50] <= data_col105[49];
   data_col105[51] <= data_col105[50];
   data_col105[52] <= data_col105[51];
   data_col105[53] <= data_col105[52];
   data_col105[54] <= data_col105[53];
   data_col105[55] <= data_col105[54];
   data_col105[56] <= data_col105[55];
   data_col105[57] <= data_col105[56];
   data_col105[58] <= data_col105[57];
   data_col105[59] <= data_col105[58];
   data_col105[60] <= data_col105[59];
   data_col105[61] <= data_col105[60];
   data_col105[62] <= data_col105[61];
   data_col105[63] <= data_col105[62];
   data_col105[64] <= data_col105[63];
   data_col105[65] <= data_col105[64];
   data_col105[66] <= data_col105[65];
   data_col105[67] <= data_col105[66];
   data_col105[68] <= data_col105[67];
   data_col105[69] <= data_col105[68];
   data_col105[70] <= data_col105[69];
   data_col105[71] <= data_col105[70];
   data_col105[72] <= data_col105[71];
   data_col105[73] <= data_col105[72];
   data_col105[74] <= data_col105[73];
   data_col105[75] <= data_col105[74];
   data_col105[76] <= data_col105[75];
   data_col105[77] <= data_col105[76];
   data_col105[78] <= data_col105[77];
   data_col105[79] <= data_col105[78];
   data_col105[80] <= data_col105[79];
   data_col105[81] <= data_col105[80];
   data_col105[82] <= data_col105[81];
   data_col105[83] <= data_col105[82];
   data_col105[84] <= data_col105[83];
   data_col105[85] <= data_col105[84];
   data_col105[86] <= data_col105[85];
   data_col105[87] <= data_col105[86];
   data_col105[88] <= data_col105[87];
   data_col105[89] <= data_col105[88];
   data_col105[90] <= data_col105[89];
   data_col105[91] <= data_col105[90];
   data_col105[92] <= data_col105[91];
   data_col105[93] <= data_col105[92];
   data_col105[94] <= data_col105[93];
   data_col105[95] <= data_col105[94];
   data_col105[96] <= data_col105[95];
   data_col105[97] <= data_col105[96];
   data_col105[98] <= data_col105[97];
   data_col105[99] <= data_col105[98];
   data_col105[100] <= data_col105[99];
   data_col105[101] <= data_col105[100];
   data_col105[102] <= data_col105[101];
   data_col105[103] <= data_col105[102];
   data_col105[104] <= data_col105[103];
   data_col105[105] <= data_col105[104];

   data_col106[1] <= data[59];
   data_col106[2] <= data_col106[1];
   data_col106[3] <= data_col106[2];
   data_col106[4] <= data_col106[3];
   data_col106[5] <= data_col106[4];
   data_col106[6] <= data_col106[5];
   data_col106[7] <= data_col106[6];
   data_col106[8] <= data_col106[7];
   data_col106[9] <= data_col106[8];
   data_col106[10] <= data_col106[9];
   data_col106[11] <= data_col106[10];
   data_col106[12] <= data_col106[11];
   data_col106[13] <= data_col106[12];
   data_col106[14] <= data_col106[13];
   data_col106[15] <= data_col106[14];
   data_col106[16] <= data_col106[15];
   data_col106[17] <= data_col106[16];
   data_col106[18] <= data_col106[17];
   data_col106[19] <= data_col106[18];
   data_col106[20] <= data_col106[19];
   data_col106[21] <= data_col106[20];
   data_col106[22] <= data_col106[21];
   data_col106[23] <= data_col106[22];
   data_col106[24] <= data_col106[23];
   data_col106[25] <= data_col106[24];
   data_col106[26] <= data_col106[25];
   data_col106[27] <= data_col106[26];
   data_col106[28] <= data_col106[27];
   data_col106[29] <= data_col106[28];
   data_col106[30] <= data_col106[29];
   data_col106[31] <= data_col106[30];
   data_col106[32] <= data_col106[31];
   data_col106[33] <= data_col106[32];
   data_col106[34] <= data_col106[33];
   data_col106[35] <= data_col106[34];
   data_col106[36] <= data_col106[35];
   data_col106[37] <= data_col106[36];
   data_col106[38] <= data_col106[37];
   data_col106[39] <= data_col106[38];
   data_col106[40] <= data_col106[39];
   data_col106[41] <= data_col106[40];
   data_col106[42] <= data_col106[41];
   data_col106[43] <= data_col106[42];
   data_col106[44] <= data_col106[43];
   data_col106[45] <= data_col106[44];
   data_col106[46] <= data_col106[45];
   data_col106[47] <= data_col106[46];
   data_col106[48] <= data_col106[47];
   data_col106[49] <= data_col106[48];
   data_col106[50] <= data_col106[49];
   data_col106[51] <= data_col106[50];
   data_col106[52] <= data_col106[51];
   data_col106[53] <= data_col106[52];
   data_col106[54] <= data_col106[53];
   data_col106[55] <= data_col106[54];
   data_col106[56] <= data_col106[55];
   data_col106[57] <= data_col106[56];
   data_col106[58] <= data_col106[57];
   data_col106[59] <= data_col106[58];
   data_col106[60] <= data_col106[59];
   data_col106[61] <= data_col106[60];
   data_col106[62] <= data_col106[61];
   data_col106[63] <= data_col106[62];
   data_col106[64] <= data_col106[63];
   data_col106[65] <= data_col106[64];
   data_col106[66] <= data_col106[65];
   data_col106[67] <= data_col106[66];
   data_col106[68] <= data_col106[67];
   data_col106[69] <= data_col106[68];
   data_col106[70] <= data_col106[69];
   data_col106[71] <= data_col106[70];
   data_col106[72] <= data_col106[71];
   data_col106[73] <= data_col106[72];
   data_col106[74] <= data_col106[73];
   data_col106[75] <= data_col106[74];
   data_col106[76] <= data_col106[75];
   data_col106[77] <= data_col106[76];
   data_col106[78] <= data_col106[77];
   data_col106[79] <= data_col106[78];
   data_col106[80] <= data_col106[79];
   data_col106[81] <= data_col106[80];
   data_col106[82] <= data_col106[81];
   data_col106[83] <= data_col106[82];
   data_col106[84] <= data_col106[83];
   data_col106[85] <= data_col106[84];
   data_col106[86] <= data_col106[85];
   data_col106[87] <= data_col106[86];
   data_col106[88] <= data_col106[87];
   data_col106[89] <= data_col106[88];
   data_col106[90] <= data_col106[89];
   data_col106[91] <= data_col106[90];
   data_col106[92] <= data_col106[91];
   data_col106[93] <= data_col106[92];
   data_col106[94] <= data_col106[93];
   data_col106[95] <= data_col106[94];
   data_col106[96] <= data_col106[95];
   data_col106[97] <= data_col106[96];
   data_col106[98] <= data_col106[97];
   data_col106[99] <= data_col106[98];
   data_col106[100] <= data_col106[99];
   data_col106[101] <= data_col106[100];
   data_col106[102] <= data_col106[101];
   data_col106[103] <= data_col106[102];
   data_col106[104] <= data_col106[103];
   data_col106[105] <= data_col106[104];
   data_col106[106] <= data_col106[105];

   data_col107[1] <= data[58];
   data_col107[2] <= data_col107[1];
   data_col107[3] <= data_col107[2];
   data_col107[4] <= data_col107[3];
   data_col107[5] <= data_col107[4];
   data_col107[6] <= data_col107[5];
   data_col107[7] <= data_col107[6];
   data_col107[8] <= data_col107[7];
   data_col107[9] <= data_col107[8];
   data_col107[10] <= data_col107[9];
   data_col107[11] <= data_col107[10];
   data_col107[12] <= data_col107[11];
   data_col107[13] <= data_col107[12];
   data_col107[14] <= data_col107[13];
   data_col107[15] <= data_col107[14];
   data_col107[16] <= data_col107[15];
   data_col107[17] <= data_col107[16];
   data_col107[18] <= data_col107[17];
   data_col107[19] <= data_col107[18];
   data_col107[20] <= data_col107[19];
   data_col107[21] <= data_col107[20];
   data_col107[22] <= data_col107[21];
   data_col107[23] <= data_col107[22];
   data_col107[24] <= data_col107[23];
   data_col107[25] <= data_col107[24];
   data_col107[26] <= data_col107[25];
   data_col107[27] <= data_col107[26];
   data_col107[28] <= data_col107[27];
   data_col107[29] <= data_col107[28];
   data_col107[30] <= data_col107[29];
   data_col107[31] <= data_col107[30];
   data_col107[32] <= data_col107[31];
   data_col107[33] <= data_col107[32];
   data_col107[34] <= data_col107[33];
   data_col107[35] <= data_col107[34];
   data_col107[36] <= data_col107[35];
   data_col107[37] <= data_col107[36];
   data_col107[38] <= data_col107[37];
   data_col107[39] <= data_col107[38];
   data_col107[40] <= data_col107[39];
   data_col107[41] <= data_col107[40];
   data_col107[42] <= data_col107[41];
   data_col107[43] <= data_col107[42];
   data_col107[44] <= data_col107[43];
   data_col107[45] <= data_col107[44];
   data_col107[46] <= data_col107[45];
   data_col107[47] <= data_col107[46];
   data_col107[48] <= data_col107[47];
   data_col107[49] <= data_col107[48];
   data_col107[50] <= data_col107[49];
   data_col107[51] <= data_col107[50];
   data_col107[52] <= data_col107[51];
   data_col107[53] <= data_col107[52];
   data_col107[54] <= data_col107[53];
   data_col107[55] <= data_col107[54];
   data_col107[56] <= data_col107[55];
   data_col107[57] <= data_col107[56];
   data_col107[58] <= data_col107[57];
   data_col107[59] <= data_col107[58];
   data_col107[60] <= data_col107[59];
   data_col107[61] <= data_col107[60];
   data_col107[62] <= data_col107[61];
   data_col107[63] <= data_col107[62];
   data_col107[64] <= data_col107[63];
   data_col107[65] <= data_col107[64];
   data_col107[66] <= data_col107[65];
   data_col107[67] <= data_col107[66];
   data_col107[68] <= data_col107[67];
   data_col107[69] <= data_col107[68];
   data_col107[70] <= data_col107[69];
   data_col107[71] <= data_col107[70];
   data_col107[72] <= data_col107[71];
   data_col107[73] <= data_col107[72];
   data_col107[74] <= data_col107[73];
   data_col107[75] <= data_col107[74];
   data_col107[76] <= data_col107[75];
   data_col107[77] <= data_col107[76];
   data_col107[78] <= data_col107[77];
   data_col107[79] <= data_col107[78];
   data_col107[80] <= data_col107[79];
   data_col107[81] <= data_col107[80];
   data_col107[82] <= data_col107[81];
   data_col107[83] <= data_col107[82];
   data_col107[84] <= data_col107[83];
   data_col107[85] <= data_col107[84];
   data_col107[86] <= data_col107[85];
   data_col107[87] <= data_col107[86];
   data_col107[88] <= data_col107[87];
   data_col107[89] <= data_col107[88];
   data_col107[90] <= data_col107[89];
   data_col107[91] <= data_col107[90];
   data_col107[92] <= data_col107[91];
   data_col107[93] <= data_col107[92];
   data_col107[94] <= data_col107[93];
   data_col107[95] <= data_col107[94];
   data_col107[96] <= data_col107[95];
   data_col107[97] <= data_col107[96];
   data_col107[98] <= data_col107[97];
   data_col107[99] <= data_col107[98];
   data_col107[100] <= data_col107[99];
   data_col107[101] <= data_col107[100];
   data_col107[102] <= data_col107[101];
   data_col107[103] <= data_col107[102];
   data_col107[104] <= data_col107[103];
   data_col107[105] <= data_col107[104];
   data_col107[106] <= data_col107[105];
   data_col107[107] <= data_col107[106];

   data_col108[1] <= data[57];
   data_col108[2] <= data_col108[1];
   data_col108[3] <= data_col108[2];
   data_col108[4] <= data_col108[3];
   data_col108[5] <= data_col108[4];
   data_col108[6] <= data_col108[5];
   data_col108[7] <= data_col108[6];
   data_col108[8] <= data_col108[7];
   data_col108[9] <= data_col108[8];
   data_col108[10] <= data_col108[9];
   data_col108[11] <= data_col108[10];
   data_col108[12] <= data_col108[11];
   data_col108[13] <= data_col108[12];
   data_col108[14] <= data_col108[13];
   data_col108[15] <= data_col108[14];
   data_col108[16] <= data_col108[15];
   data_col108[17] <= data_col108[16];
   data_col108[18] <= data_col108[17];
   data_col108[19] <= data_col108[18];
   data_col108[20] <= data_col108[19];
   data_col108[21] <= data_col108[20];
   data_col108[22] <= data_col108[21];
   data_col108[23] <= data_col108[22];
   data_col108[24] <= data_col108[23];
   data_col108[25] <= data_col108[24];
   data_col108[26] <= data_col108[25];
   data_col108[27] <= data_col108[26];
   data_col108[28] <= data_col108[27];
   data_col108[29] <= data_col108[28];
   data_col108[30] <= data_col108[29];
   data_col108[31] <= data_col108[30];
   data_col108[32] <= data_col108[31];
   data_col108[33] <= data_col108[32];
   data_col108[34] <= data_col108[33];
   data_col108[35] <= data_col108[34];
   data_col108[36] <= data_col108[35];
   data_col108[37] <= data_col108[36];
   data_col108[38] <= data_col108[37];
   data_col108[39] <= data_col108[38];
   data_col108[40] <= data_col108[39];
   data_col108[41] <= data_col108[40];
   data_col108[42] <= data_col108[41];
   data_col108[43] <= data_col108[42];
   data_col108[44] <= data_col108[43];
   data_col108[45] <= data_col108[44];
   data_col108[46] <= data_col108[45];
   data_col108[47] <= data_col108[46];
   data_col108[48] <= data_col108[47];
   data_col108[49] <= data_col108[48];
   data_col108[50] <= data_col108[49];
   data_col108[51] <= data_col108[50];
   data_col108[52] <= data_col108[51];
   data_col108[53] <= data_col108[52];
   data_col108[54] <= data_col108[53];
   data_col108[55] <= data_col108[54];
   data_col108[56] <= data_col108[55];
   data_col108[57] <= data_col108[56];
   data_col108[58] <= data_col108[57];
   data_col108[59] <= data_col108[58];
   data_col108[60] <= data_col108[59];
   data_col108[61] <= data_col108[60];
   data_col108[62] <= data_col108[61];
   data_col108[63] <= data_col108[62];
   data_col108[64] <= data_col108[63];
   data_col108[65] <= data_col108[64];
   data_col108[66] <= data_col108[65];
   data_col108[67] <= data_col108[66];
   data_col108[68] <= data_col108[67];
   data_col108[69] <= data_col108[68];
   data_col108[70] <= data_col108[69];
   data_col108[71] <= data_col108[70];
   data_col108[72] <= data_col108[71];
   data_col108[73] <= data_col108[72];
   data_col108[74] <= data_col108[73];
   data_col108[75] <= data_col108[74];
   data_col108[76] <= data_col108[75];
   data_col108[77] <= data_col108[76];
   data_col108[78] <= data_col108[77];
   data_col108[79] <= data_col108[78];
   data_col108[80] <= data_col108[79];
   data_col108[81] <= data_col108[80];
   data_col108[82] <= data_col108[81];
   data_col108[83] <= data_col108[82];
   data_col108[84] <= data_col108[83];
   data_col108[85] <= data_col108[84];
   data_col108[86] <= data_col108[85];
   data_col108[87] <= data_col108[86];
   data_col108[88] <= data_col108[87];
   data_col108[89] <= data_col108[88];
   data_col108[90] <= data_col108[89];
   data_col108[91] <= data_col108[90];
   data_col108[92] <= data_col108[91];
   data_col108[93] <= data_col108[92];
   data_col108[94] <= data_col108[93];
   data_col108[95] <= data_col108[94];
   data_col108[96] <= data_col108[95];
   data_col108[97] <= data_col108[96];
   data_col108[98] <= data_col108[97];
   data_col108[99] <= data_col108[98];
   data_col108[100] <= data_col108[99];
   data_col108[101] <= data_col108[100];
   data_col108[102] <= data_col108[101];
   data_col108[103] <= data_col108[102];
   data_col108[104] <= data_col108[103];
   data_col108[105] <= data_col108[104];
   data_col108[106] <= data_col108[105];
   data_col108[107] <= data_col108[106];
   data_col108[108] <= data_col108[107];

   data_col109[1] <= data[56];
   data_col109[2] <= data_col109[1];
   data_col109[3] <= data_col109[2];
   data_col109[4] <= data_col109[3];
   data_col109[5] <= data_col109[4];
   data_col109[6] <= data_col109[5];
   data_col109[7] <= data_col109[6];
   data_col109[8] <= data_col109[7];
   data_col109[9] <= data_col109[8];
   data_col109[10] <= data_col109[9];
   data_col109[11] <= data_col109[10];
   data_col109[12] <= data_col109[11];
   data_col109[13] <= data_col109[12];
   data_col109[14] <= data_col109[13];
   data_col109[15] <= data_col109[14];
   data_col109[16] <= data_col109[15];
   data_col109[17] <= data_col109[16];
   data_col109[18] <= data_col109[17];
   data_col109[19] <= data_col109[18];
   data_col109[20] <= data_col109[19];
   data_col109[21] <= data_col109[20];
   data_col109[22] <= data_col109[21];
   data_col109[23] <= data_col109[22];
   data_col109[24] <= data_col109[23];
   data_col109[25] <= data_col109[24];
   data_col109[26] <= data_col109[25];
   data_col109[27] <= data_col109[26];
   data_col109[28] <= data_col109[27];
   data_col109[29] <= data_col109[28];
   data_col109[30] <= data_col109[29];
   data_col109[31] <= data_col109[30];
   data_col109[32] <= data_col109[31];
   data_col109[33] <= data_col109[32];
   data_col109[34] <= data_col109[33];
   data_col109[35] <= data_col109[34];
   data_col109[36] <= data_col109[35];
   data_col109[37] <= data_col109[36];
   data_col109[38] <= data_col109[37];
   data_col109[39] <= data_col109[38];
   data_col109[40] <= data_col109[39];
   data_col109[41] <= data_col109[40];
   data_col109[42] <= data_col109[41];
   data_col109[43] <= data_col109[42];
   data_col109[44] <= data_col109[43];
   data_col109[45] <= data_col109[44];
   data_col109[46] <= data_col109[45];
   data_col109[47] <= data_col109[46];
   data_col109[48] <= data_col109[47];
   data_col109[49] <= data_col109[48];
   data_col109[50] <= data_col109[49];
   data_col109[51] <= data_col109[50];
   data_col109[52] <= data_col109[51];
   data_col109[53] <= data_col109[52];
   data_col109[54] <= data_col109[53];
   data_col109[55] <= data_col109[54];
   data_col109[56] <= data_col109[55];
   data_col109[57] <= data_col109[56];
   data_col109[58] <= data_col109[57];
   data_col109[59] <= data_col109[58];
   data_col109[60] <= data_col109[59];
   data_col109[61] <= data_col109[60];
   data_col109[62] <= data_col109[61];
   data_col109[63] <= data_col109[62];
   data_col109[64] <= data_col109[63];
   data_col109[65] <= data_col109[64];
   data_col109[66] <= data_col109[65];
   data_col109[67] <= data_col109[66];
   data_col109[68] <= data_col109[67];
   data_col109[69] <= data_col109[68];
   data_col109[70] <= data_col109[69];
   data_col109[71] <= data_col109[70];
   data_col109[72] <= data_col109[71];
   data_col109[73] <= data_col109[72];
   data_col109[74] <= data_col109[73];
   data_col109[75] <= data_col109[74];
   data_col109[76] <= data_col109[75];
   data_col109[77] <= data_col109[76];
   data_col109[78] <= data_col109[77];
   data_col109[79] <= data_col109[78];
   data_col109[80] <= data_col109[79];
   data_col109[81] <= data_col109[80];
   data_col109[82] <= data_col109[81];
   data_col109[83] <= data_col109[82];
   data_col109[84] <= data_col109[83];
   data_col109[85] <= data_col109[84];
   data_col109[86] <= data_col109[85];
   data_col109[87] <= data_col109[86];
   data_col109[88] <= data_col109[87];
   data_col109[89] <= data_col109[88];
   data_col109[90] <= data_col109[89];
   data_col109[91] <= data_col109[90];
   data_col109[92] <= data_col109[91];
   data_col109[93] <= data_col109[92];
   data_col109[94] <= data_col109[93];
   data_col109[95] <= data_col109[94];
   data_col109[96] <= data_col109[95];
   data_col109[97] <= data_col109[96];
   data_col109[98] <= data_col109[97];
   data_col109[99] <= data_col109[98];
   data_col109[100] <= data_col109[99];
   data_col109[101] <= data_col109[100];
   data_col109[102] <= data_col109[101];
   data_col109[103] <= data_col109[102];
   data_col109[104] <= data_col109[103];
   data_col109[105] <= data_col109[104];
   data_col109[106] <= data_col109[105];
   data_col109[107] <= data_col109[106];
   data_col109[108] <= data_col109[107];
   data_col109[109] <= data_col109[108];

   data_col110[1] <= data[55];
   data_col110[2] <= data_col110[1];
   data_col110[3] <= data_col110[2];
   data_col110[4] <= data_col110[3];
   data_col110[5] <= data_col110[4];
   data_col110[6] <= data_col110[5];
   data_col110[7] <= data_col110[6];
   data_col110[8] <= data_col110[7];
   data_col110[9] <= data_col110[8];
   data_col110[10] <= data_col110[9];
   data_col110[11] <= data_col110[10];
   data_col110[12] <= data_col110[11];
   data_col110[13] <= data_col110[12];
   data_col110[14] <= data_col110[13];
   data_col110[15] <= data_col110[14];
   data_col110[16] <= data_col110[15];
   data_col110[17] <= data_col110[16];
   data_col110[18] <= data_col110[17];
   data_col110[19] <= data_col110[18];
   data_col110[20] <= data_col110[19];
   data_col110[21] <= data_col110[20];
   data_col110[22] <= data_col110[21];
   data_col110[23] <= data_col110[22];
   data_col110[24] <= data_col110[23];
   data_col110[25] <= data_col110[24];
   data_col110[26] <= data_col110[25];
   data_col110[27] <= data_col110[26];
   data_col110[28] <= data_col110[27];
   data_col110[29] <= data_col110[28];
   data_col110[30] <= data_col110[29];
   data_col110[31] <= data_col110[30];
   data_col110[32] <= data_col110[31];
   data_col110[33] <= data_col110[32];
   data_col110[34] <= data_col110[33];
   data_col110[35] <= data_col110[34];
   data_col110[36] <= data_col110[35];
   data_col110[37] <= data_col110[36];
   data_col110[38] <= data_col110[37];
   data_col110[39] <= data_col110[38];
   data_col110[40] <= data_col110[39];
   data_col110[41] <= data_col110[40];
   data_col110[42] <= data_col110[41];
   data_col110[43] <= data_col110[42];
   data_col110[44] <= data_col110[43];
   data_col110[45] <= data_col110[44];
   data_col110[46] <= data_col110[45];
   data_col110[47] <= data_col110[46];
   data_col110[48] <= data_col110[47];
   data_col110[49] <= data_col110[48];
   data_col110[50] <= data_col110[49];
   data_col110[51] <= data_col110[50];
   data_col110[52] <= data_col110[51];
   data_col110[53] <= data_col110[52];
   data_col110[54] <= data_col110[53];
   data_col110[55] <= data_col110[54];
   data_col110[56] <= data_col110[55];
   data_col110[57] <= data_col110[56];
   data_col110[58] <= data_col110[57];
   data_col110[59] <= data_col110[58];
   data_col110[60] <= data_col110[59];
   data_col110[61] <= data_col110[60];
   data_col110[62] <= data_col110[61];
   data_col110[63] <= data_col110[62];
   data_col110[64] <= data_col110[63];
   data_col110[65] <= data_col110[64];
   data_col110[66] <= data_col110[65];
   data_col110[67] <= data_col110[66];
   data_col110[68] <= data_col110[67];
   data_col110[69] <= data_col110[68];
   data_col110[70] <= data_col110[69];
   data_col110[71] <= data_col110[70];
   data_col110[72] <= data_col110[71];
   data_col110[73] <= data_col110[72];
   data_col110[74] <= data_col110[73];
   data_col110[75] <= data_col110[74];
   data_col110[76] <= data_col110[75];
   data_col110[77] <= data_col110[76];
   data_col110[78] <= data_col110[77];
   data_col110[79] <= data_col110[78];
   data_col110[80] <= data_col110[79];
   data_col110[81] <= data_col110[80];
   data_col110[82] <= data_col110[81];
   data_col110[83] <= data_col110[82];
   data_col110[84] <= data_col110[83];
   data_col110[85] <= data_col110[84];
   data_col110[86] <= data_col110[85];
   data_col110[87] <= data_col110[86];
   data_col110[88] <= data_col110[87];
   data_col110[89] <= data_col110[88];
   data_col110[90] <= data_col110[89];
   data_col110[91] <= data_col110[90];
   data_col110[92] <= data_col110[91];
   data_col110[93] <= data_col110[92];
   data_col110[94] <= data_col110[93];
   data_col110[95] <= data_col110[94];
   data_col110[96] <= data_col110[95];
   data_col110[97] <= data_col110[96];
   data_col110[98] <= data_col110[97];
   data_col110[99] <= data_col110[98];
   data_col110[100] <= data_col110[99];
   data_col110[101] <= data_col110[100];
   data_col110[102] <= data_col110[101];
   data_col110[103] <= data_col110[102];
   data_col110[104] <= data_col110[103];
   data_col110[105] <= data_col110[104];
   data_col110[106] <= data_col110[105];
   data_col110[107] <= data_col110[106];
   data_col110[108] <= data_col110[107];
   data_col110[109] <= data_col110[108];
   data_col110[110] <= data_col110[109];

   data_col111[1] <= data[54];
   data_col111[2] <= data_col111[1];
   data_col111[3] <= data_col111[2];
   data_col111[4] <= data_col111[3];
   data_col111[5] <= data_col111[4];
   data_col111[6] <= data_col111[5];
   data_col111[7] <= data_col111[6];
   data_col111[8] <= data_col111[7];
   data_col111[9] <= data_col111[8];
   data_col111[10] <= data_col111[9];
   data_col111[11] <= data_col111[10];
   data_col111[12] <= data_col111[11];
   data_col111[13] <= data_col111[12];
   data_col111[14] <= data_col111[13];
   data_col111[15] <= data_col111[14];
   data_col111[16] <= data_col111[15];
   data_col111[17] <= data_col111[16];
   data_col111[18] <= data_col111[17];
   data_col111[19] <= data_col111[18];
   data_col111[20] <= data_col111[19];
   data_col111[21] <= data_col111[20];
   data_col111[22] <= data_col111[21];
   data_col111[23] <= data_col111[22];
   data_col111[24] <= data_col111[23];
   data_col111[25] <= data_col111[24];
   data_col111[26] <= data_col111[25];
   data_col111[27] <= data_col111[26];
   data_col111[28] <= data_col111[27];
   data_col111[29] <= data_col111[28];
   data_col111[30] <= data_col111[29];
   data_col111[31] <= data_col111[30];
   data_col111[32] <= data_col111[31];
   data_col111[33] <= data_col111[32];
   data_col111[34] <= data_col111[33];
   data_col111[35] <= data_col111[34];
   data_col111[36] <= data_col111[35];
   data_col111[37] <= data_col111[36];
   data_col111[38] <= data_col111[37];
   data_col111[39] <= data_col111[38];
   data_col111[40] <= data_col111[39];
   data_col111[41] <= data_col111[40];
   data_col111[42] <= data_col111[41];
   data_col111[43] <= data_col111[42];
   data_col111[44] <= data_col111[43];
   data_col111[45] <= data_col111[44];
   data_col111[46] <= data_col111[45];
   data_col111[47] <= data_col111[46];
   data_col111[48] <= data_col111[47];
   data_col111[49] <= data_col111[48];
   data_col111[50] <= data_col111[49];
   data_col111[51] <= data_col111[50];
   data_col111[52] <= data_col111[51];
   data_col111[53] <= data_col111[52];
   data_col111[54] <= data_col111[53];
   data_col111[55] <= data_col111[54];
   data_col111[56] <= data_col111[55];
   data_col111[57] <= data_col111[56];
   data_col111[58] <= data_col111[57];
   data_col111[59] <= data_col111[58];
   data_col111[60] <= data_col111[59];
   data_col111[61] <= data_col111[60];
   data_col111[62] <= data_col111[61];
   data_col111[63] <= data_col111[62];
   data_col111[64] <= data_col111[63];
   data_col111[65] <= data_col111[64];
   data_col111[66] <= data_col111[65];
   data_col111[67] <= data_col111[66];
   data_col111[68] <= data_col111[67];
   data_col111[69] <= data_col111[68];
   data_col111[70] <= data_col111[69];
   data_col111[71] <= data_col111[70];
   data_col111[72] <= data_col111[71];
   data_col111[73] <= data_col111[72];
   data_col111[74] <= data_col111[73];
   data_col111[75] <= data_col111[74];
   data_col111[76] <= data_col111[75];
   data_col111[77] <= data_col111[76];
   data_col111[78] <= data_col111[77];
   data_col111[79] <= data_col111[78];
   data_col111[80] <= data_col111[79];
   data_col111[81] <= data_col111[80];
   data_col111[82] <= data_col111[81];
   data_col111[83] <= data_col111[82];
   data_col111[84] <= data_col111[83];
   data_col111[85] <= data_col111[84];
   data_col111[86] <= data_col111[85];
   data_col111[87] <= data_col111[86];
   data_col111[88] <= data_col111[87];
   data_col111[89] <= data_col111[88];
   data_col111[90] <= data_col111[89];
   data_col111[91] <= data_col111[90];
   data_col111[92] <= data_col111[91];
   data_col111[93] <= data_col111[92];
   data_col111[94] <= data_col111[93];
   data_col111[95] <= data_col111[94];
   data_col111[96] <= data_col111[95];
   data_col111[97] <= data_col111[96];
   data_col111[98] <= data_col111[97];
   data_col111[99] <= data_col111[98];
   data_col111[100] <= data_col111[99];
   data_col111[101] <= data_col111[100];
   data_col111[102] <= data_col111[101];
   data_col111[103] <= data_col111[102];
   data_col111[104] <= data_col111[103];
   data_col111[105] <= data_col111[104];
   data_col111[106] <= data_col111[105];
   data_col111[107] <= data_col111[106];
   data_col111[108] <= data_col111[107];
   data_col111[109] <= data_col111[108];
   data_col111[110] <= data_col111[109];
   data_col111[111] <= data_col111[110];

   data_col112[1] <= data[53];
   data_col112[2] <= data_col112[1];
   data_col112[3] <= data_col112[2];
   data_col112[4] <= data_col112[3];
   data_col112[5] <= data_col112[4];
   data_col112[6] <= data_col112[5];
   data_col112[7] <= data_col112[6];
   data_col112[8] <= data_col112[7];
   data_col112[9] <= data_col112[8];
   data_col112[10] <= data_col112[9];
   data_col112[11] <= data_col112[10];
   data_col112[12] <= data_col112[11];
   data_col112[13] <= data_col112[12];
   data_col112[14] <= data_col112[13];
   data_col112[15] <= data_col112[14];
   data_col112[16] <= data_col112[15];
   data_col112[17] <= data_col112[16];
   data_col112[18] <= data_col112[17];
   data_col112[19] <= data_col112[18];
   data_col112[20] <= data_col112[19];
   data_col112[21] <= data_col112[20];
   data_col112[22] <= data_col112[21];
   data_col112[23] <= data_col112[22];
   data_col112[24] <= data_col112[23];
   data_col112[25] <= data_col112[24];
   data_col112[26] <= data_col112[25];
   data_col112[27] <= data_col112[26];
   data_col112[28] <= data_col112[27];
   data_col112[29] <= data_col112[28];
   data_col112[30] <= data_col112[29];
   data_col112[31] <= data_col112[30];
   data_col112[32] <= data_col112[31];
   data_col112[33] <= data_col112[32];
   data_col112[34] <= data_col112[33];
   data_col112[35] <= data_col112[34];
   data_col112[36] <= data_col112[35];
   data_col112[37] <= data_col112[36];
   data_col112[38] <= data_col112[37];
   data_col112[39] <= data_col112[38];
   data_col112[40] <= data_col112[39];
   data_col112[41] <= data_col112[40];
   data_col112[42] <= data_col112[41];
   data_col112[43] <= data_col112[42];
   data_col112[44] <= data_col112[43];
   data_col112[45] <= data_col112[44];
   data_col112[46] <= data_col112[45];
   data_col112[47] <= data_col112[46];
   data_col112[48] <= data_col112[47];
   data_col112[49] <= data_col112[48];
   data_col112[50] <= data_col112[49];
   data_col112[51] <= data_col112[50];
   data_col112[52] <= data_col112[51];
   data_col112[53] <= data_col112[52];
   data_col112[54] <= data_col112[53];
   data_col112[55] <= data_col112[54];
   data_col112[56] <= data_col112[55];
   data_col112[57] <= data_col112[56];
   data_col112[58] <= data_col112[57];
   data_col112[59] <= data_col112[58];
   data_col112[60] <= data_col112[59];
   data_col112[61] <= data_col112[60];
   data_col112[62] <= data_col112[61];
   data_col112[63] <= data_col112[62];
   data_col112[64] <= data_col112[63];
   data_col112[65] <= data_col112[64];
   data_col112[66] <= data_col112[65];
   data_col112[67] <= data_col112[66];
   data_col112[68] <= data_col112[67];
   data_col112[69] <= data_col112[68];
   data_col112[70] <= data_col112[69];
   data_col112[71] <= data_col112[70];
   data_col112[72] <= data_col112[71];
   data_col112[73] <= data_col112[72];
   data_col112[74] <= data_col112[73];
   data_col112[75] <= data_col112[74];
   data_col112[76] <= data_col112[75];
   data_col112[77] <= data_col112[76];
   data_col112[78] <= data_col112[77];
   data_col112[79] <= data_col112[78];
   data_col112[80] <= data_col112[79];
   data_col112[81] <= data_col112[80];
   data_col112[82] <= data_col112[81];
   data_col112[83] <= data_col112[82];
   data_col112[84] <= data_col112[83];
   data_col112[85] <= data_col112[84];
   data_col112[86] <= data_col112[85];
   data_col112[87] <= data_col112[86];
   data_col112[88] <= data_col112[87];
   data_col112[89] <= data_col112[88];
   data_col112[90] <= data_col112[89];
   data_col112[91] <= data_col112[90];
   data_col112[92] <= data_col112[91];
   data_col112[93] <= data_col112[92];
   data_col112[94] <= data_col112[93];
   data_col112[95] <= data_col112[94];
   data_col112[96] <= data_col112[95];
   data_col112[97] <= data_col112[96];
   data_col112[98] <= data_col112[97];
   data_col112[99] <= data_col112[98];
   data_col112[100] <= data_col112[99];
   data_col112[101] <= data_col112[100];
   data_col112[102] <= data_col112[101];
   data_col112[103] <= data_col112[102];
   data_col112[104] <= data_col112[103];
   data_col112[105] <= data_col112[104];
   data_col112[106] <= data_col112[105];
   data_col112[107] <= data_col112[106];
   data_col112[108] <= data_col112[107];
   data_col112[109] <= data_col112[108];
   data_col112[110] <= data_col112[109];
   data_col112[111] <= data_col112[110];
   data_col112[112] <= data_col112[111];

   data_col113[1] <= data[52];
   data_col113[2] <= data_col113[1];
   data_col113[3] <= data_col113[2];
   data_col113[4] <= data_col113[3];
   data_col113[5] <= data_col113[4];
   data_col113[6] <= data_col113[5];
   data_col113[7] <= data_col113[6];
   data_col113[8] <= data_col113[7];
   data_col113[9] <= data_col113[8];
   data_col113[10] <= data_col113[9];
   data_col113[11] <= data_col113[10];
   data_col113[12] <= data_col113[11];
   data_col113[13] <= data_col113[12];
   data_col113[14] <= data_col113[13];
   data_col113[15] <= data_col113[14];
   data_col113[16] <= data_col113[15];
   data_col113[17] <= data_col113[16];
   data_col113[18] <= data_col113[17];
   data_col113[19] <= data_col113[18];
   data_col113[20] <= data_col113[19];
   data_col113[21] <= data_col113[20];
   data_col113[22] <= data_col113[21];
   data_col113[23] <= data_col113[22];
   data_col113[24] <= data_col113[23];
   data_col113[25] <= data_col113[24];
   data_col113[26] <= data_col113[25];
   data_col113[27] <= data_col113[26];
   data_col113[28] <= data_col113[27];
   data_col113[29] <= data_col113[28];
   data_col113[30] <= data_col113[29];
   data_col113[31] <= data_col113[30];
   data_col113[32] <= data_col113[31];
   data_col113[33] <= data_col113[32];
   data_col113[34] <= data_col113[33];
   data_col113[35] <= data_col113[34];
   data_col113[36] <= data_col113[35];
   data_col113[37] <= data_col113[36];
   data_col113[38] <= data_col113[37];
   data_col113[39] <= data_col113[38];
   data_col113[40] <= data_col113[39];
   data_col113[41] <= data_col113[40];
   data_col113[42] <= data_col113[41];
   data_col113[43] <= data_col113[42];
   data_col113[44] <= data_col113[43];
   data_col113[45] <= data_col113[44];
   data_col113[46] <= data_col113[45];
   data_col113[47] <= data_col113[46];
   data_col113[48] <= data_col113[47];
   data_col113[49] <= data_col113[48];
   data_col113[50] <= data_col113[49];
   data_col113[51] <= data_col113[50];
   data_col113[52] <= data_col113[51];
   data_col113[53] <= data_col113[52];
   data_col113[54] <= data_col113[53];
   data_col113[55] <= data_col113[54];
   data_col113[56] <= data_col113[55];
   data_col113[57] <= data_col113[56];
   data_col113[58] <= data_col113[57];
   data_col113[59] <= data_col113[58];
   data_col113[60] <= data_col113[59];
   data_col113[61] <= data_col113[60];
   data_col113[62] <= data_col113[61];
   data_col113[63] <= data_col113[62];
   data_col113[64] <= data_col113[63];
   data_col113[65] <= data_col113[64];
   data_col113[66] <= data_col113[65];
   data_col113[67] <= data_col113[66];
   data_col113[68] <= data_col113[67];
   data_col113[69] <= data_col113[68];
   data_col113[70] <= data_col113[69];
   data_col113[71] <= data_col113[70];
   data_col113[72] <= data_col113[71];
   data_col113[73] <= data_col113[72];
   data_col113[74] <= data_col113[73];
   data_col113[75] <= data_col113[74];
   data_col113[76] <= data_col113[75];
   data_col113[77] <= data_col113[76];
   data_col113[78] <= data_col113[77];
   data_col113[79] <= data_col113[78];
   data_col113[80] <= data_col113[79];
   data_col113[81] <= data_col113[80];
   data_col113[82] <= data_col113[81];
   data_col113[83] <= data_col113[82];
   data_col113[84] <= data_col113[83];
   data_col113[85] <= data_col113[84];
   data_col113[86] <= data_col113[85];
   data_col113[87] <= data_col113[86];
   data_col113[88] <= data_col113[87];
   data_col113[89] <= data_col113[88];
   data_col113[90] <= data_col113[89];
   data_col113[91] <= data_col113[90];
   data_col113[92] <= data_col113[91];
   data_col113[93] <= data_col113[92];
   data_col113[94] <= data_col113[93];
   data_col113[95] <= data_col113[94];
   data_col113[96] <= data_col113[95];
   data_col113[97] <= data_col113[96];
   data_col113[98] <= data_col113[97];
   data_col113[99] <= data_col113[98];
   data_col113[100] <= data_col113[99];
   data_col113[101] <= data_col113[100];
   data_col113[102] <= data_col113[101];
   data_col113[103] <= data_col113[102];
   data_col113[104] <= data_col113[103];
   data_col113[105] <= data_col113[104];
   data_col113[106] <= data_col113[105];
   data_col113[107] <= data_col113[106];
   data_col113[108] <= data_col113[107];
   data_col113[109] <= data_col113[108];
   data_col113[110] <= data_col113[109];
   data_col113[111] <= data_col113[110];
   data_col113[112] <= data_col113[111];
   data_col113[113] <= data_col113[112];

   data_col114[1] <= data[51];
   data_col114[2] <= data_col114[1];
   data_col114[3] <= data_col114[2];
   data_col114[4] <= data_col114[3];
   data_col114[5] <= data_col114[4];
   data_col114[6] <= data_col114[5];
   data_col114[7] <= data_col114[6];
   data_col114[8] <= data_col114[7];
   data_col114[9] <= data_col114[8];
   data_col114[10] <= data_col114[9];
   data_col114[11] <= data_col114[10];
   data_col114[12] <= data_col114[11];
   data_col114[13] <= data_col114[12];
   data_col114[14] <= data_col114[13];
   data_col114[15] <= data_col114[14];
   data_col114[16] <= data_col114[15];
   data_col114[17] <= data_col114[16];
   data_col114[18] <= data_col114[17];
   data_col114[19] <= data_col114[18];
   data_col114[20] <= data_col114[19];
   data_col114[21] <= data_col114[20];
   data_col114[22] <= data_col114[21];
   data_col114[23] <= data_col114[22];
   data_col114[24] <= data_col114[23];
   data_col114[25] <= data_col114[24];
   data_col114[26] <= data_col114[25];
   data_col114[27] <= data_col114[26];
   data_col114[28] <= data_col114[27];
   data_col114[29] <= data_col114[28];
   data_col114[30] <= data_col114[29];
   data_col114[31] <= data_col114[30];
   data_col114[32] <= data_col114[31];
   data_col114[33] <= data_col114[32];
   data_col114[34] <= data_col114[33];
   data_col114[35] <= data_col114[34];
   data_col114[36] <= data_col114[35];
   data_col114[37] <= data_col114[36];
   data_col114[38] <= data_col114[37];
   data_col114[39] <= data_col114[38];
   data_col114[40] <= data_col114[39];
   data_col114[41] <= data_col114[40];
   data_col114[42] <= data_col114[41];
   data_col114[43] <= data_col114[42];
   data_col114[44] <= data_col114[43];
   data_col114[45] <= data_col114[44];
   data_col114[46] <= data_col114[45];
   data_col114[47] <= data_col114[46];
   data_col114[48] <= data_col114[47];
   data_col114[49] <= data_col114[48];
   data_col114[50] <= data_col114[49];
   data_col114[51] <= data_col114[50];
   data_col114[52] <= data_col114[51];
   data_col114[53] <= data_col114[52];
   data_col114[54] <= data_col114[53];
   data_col114[55] <= data_col114[54];
   data_col114[56] <= data_col114[55];
   data_col114[57] <= data_col114[56];
   data_col114[58] <= data_col114[57];
   data_col114[59] <= data_col114[58];
   data_col114[60] <= data_col114[59];
   data_col114[61] <= data_col114[60];
   data_col114[62] <= data_col114[61];
   data_col114[63] <= data_col114[62];
   data_col114[64] <= data_col114[63];
   data_col114[65] <= data_col114[64];
   data_col114[66] <= data_col114[65];
   data_col114[67] <= data_col114[66];
   data_col114[68] <= data_col114[67];
   data_col114[69] <= data_col114[68];
   data_col114[70] <= data_col114[69];
   data_col114[71] <= data_col114[70];
   data_col114[72] <= data_col114[71];
   data_col114[73] <= data_col114[72];
   data_col114[74] <= data_col114[73];
   data_col114[75] <= data_col114[74];
   data_col114[76] <= data_col114[75];
   data_col114[77] <= data_col114[76];
   data_col114[78] <= data_col114[77];
   data_col114[79] <= data_col114[78];
   data_col114[80] <= data_col114[79];
   data_col114[81] <= data_col114[80];
   data_col114[82] <= data_col114[81];
   data_col114[83] <= data_col114[82];
   data_col114[84] <= data_col114[83];
   data_col114[85] <= data_col114[84];
   data_col114[86] <= data_col114[85];
   data_col114[87] <= data_col114[86];
   data_col114[88] <= data_col114[87];
   data_col114[89] <= data_col114[88];
   data_col114[90] <= data_col114[89];
   data_col114[91] <= data_col114[90];
   data_col114[92] <= data_col114[91];
   data_col114[93] <= data_col114[92];
   data_col114[94] <= data_col114[93];
   data_col114[95] <= data_col114[94];
   data_col114[96] <= data_col114[95];
   data_col114[97] <= data_col114[96];
   data_col114[98] <= data_col114[97];
   data_col114[99] <= data_col114[98];
   data_col114[100] <= data_col114[99];
   data_col114[101] <= data_col114[100];
   data_col114[102] <= data_col114[101];
   data_col114[103] <= data_col114[102];
   data_col114[104] <= data_col114[103];
   data_col114[105] <= data_col114[104];
   data_col114[106] <= data_col114[105];
   data_col114[107] <= data_col114[106];
   data_col114[108] <= data_col114[107];
   data_col114[109] <= data_col114[108];
   data_col114[110] <= data_col114[109];
   data_col114[111] <= data_col114[110];
   data_col114[112] <= data_col114[111];
   data_col114[113] <= data_col114[112];
   data_col114[114] <= data_col114[113];

   data_col115[1] <= data[50];
   data_col115[2] <= data_col115[1];
   data_col115[3] <= data_col115[2];
   data_col115[4] <= data_col115[3];
   data_col115[5] <= data_col115[4];
   data_col115[6] <= data_col115[5];
   data_col115[7] <= data_col115[6];
   data_col115[8] <= data_col115[7];
   data_col115[9] <= data_col115[8];
   data_col115[10] <= data_col115[9];
   data_col115[11] <= data_col115[10];
   data_col115[12] <= data_col115[11];
   data_col115[13] <= data_col115[12];
   data_col115[14] <= data_col115[13];
   data_col115[15] <= data_col115[14];
   data_col115[16] <= data_col115[15];
   data_col115[17] <= data_col115[16];
   data_col115[18] <= data_col115[17];
   data_col115[19] <= data_col115[18];
   data_col115[20] <= data_col115[19];
   data_col115[21] <= data_col115[20];
   data_col115[22] <= data_col115[21];
   data_col115[23] <= data_col115[22];
   data_col115[24] <= data_col115[23];
   data_col115[25] <= data_col115[24];
   data_col115[26] <= data_col115[25];
   data_col115[27] <= data_col115[26];
   data_col115[28] <= data_col115[27];
   data_col115[29] <= data_col115[28];
   data_col115[30] <= data_col115[29];
   data_col115[31] <= data_col115[30];
   data_col115[32] <= data_col115[31];
   data_col115[33] <= data_col115[32];
   data_col115[34] <= data_col115[33];
   data_col115[35] <= data_col115[34];
   data_col115[36] <= data_col115[35];
   data_col115[37] <= data_col115[36];
   data_col115[38] <= data_col115[37];
   data_col115[39] <= data_col115[38];
   data_col115[40] <= data_col115[39];
   data_col115[41] <= data_col115[40];
   data_col115[42] <= data_col115[41];
   data_col115[43] <= data_col115[42];
   data_col115[44] <= data_col115[43];
   data_col115[45] <= data_col115[44];
   data_col115[46] <= data_col115[45];
   data_col115[47] <= data_col115[46];
   data_col115[48] <= data_col115[47];
   data_col115[49] <= data_col115[48];
   data_col115[50] <= data_col115[49];
   data_col115[51] <= data_col115[50];
   data_col115[52] <= data_col115[51];
   data_col115[53] <= data_col115[52];
   data_col115[54] <= data_col115[53];
   data_col115[55] <= data_col115[54];
   data_col115[56] <= data_col115[55];
   data_col115[57] <= data_col115[56];
   data_col115[58] <= data_col115[57];
   data_col115[59] <= data_col115[58];
   data_col115[60] <= data_col115[59];
   data_col115[61] <= data_col115[60];
   data_col115[62] <= data_col115[61];
   data_col115[63] <= data_col115[62];
   data_col115[64] <= data_col115[63];
   data_col115[65] <= data_col115[64];
   data_col115[66] <= data_col115[65];
   data_col115[67] <= data_col115[66];
   data_col115[68] <= data_col115[67];
   data_col115[69] <= data_col115[68];
   data_col115[70] <= data_col115[69];
   data_col115[71] <= data_col115[70];
   data_col115[72] <= data_col115[71];
   data_col115[73] <= data_col115[72];
   data_col115[74] <= data_col115[73];
   data_col115[75] <= data_col115[74];
   data_col115[76] <= data_col115[75];
   data_col115[77] <= data_col115[76];
   data_col115[78] <= data_col115[77];
   data_col115[79] <= data_col115[78];
   data_col115[80] <= data_col115[79];
   data_col115[81] <= data_col115[80];
   data_col115[82] <= data_col115[81];
   data_col115[83] <= data_col115[82];
   data_col115[84] <= data_col115[83];
   data_col115[85] <= data_col115[84];
   data_col115[86] <= data_col115[85];
   data_col115[87] <= data_col115[86];
   data_col115[88] <= data_col115[87];
   data_col115[89] <= data_col115[88];
   data_col115[90] <= data_col115[89];
   data_col115[91] <= data_col115[90];
   data_col115[92] <= data_col115[91];
   data_col115[93] <= data_col115[92];
   data_col115[94] <= data_col115[93];
   data_col115[95] <= data_col115[94];
   data_col115[96] <= data_col115[95];
   data_col115[97] <= data_col115[96];
   data_col115[98] <= data_col115[97];
   data_col115[99] <= data_col115[98];
   data_col115[100] <= data_col115[99];
   data_col115[101] <= data_col115[100];
   data_col115[102] <= data_col115[101];
   data_col115[103] <= data_col115[102];
   data_col115[104] <= data_col115[103];
   data_col115[105] <= data_col115[104];
   data_col115[106] <= data_col115[105];
   data_col115[107] <= data_col115[106];
   data_col115[108] <= data_col115[107];
   data_col115[109] <= data_col115[108];
   data_col115[110] <= data_col115[109];
   data_col115[111] <= data_col115[110];
   data_col115[112] <= data_col115[111];
   data_col115[113] <= data_col115[112];
   data_col115[114] <= data_col115[113];
   data_col115[115] <= data_col115[114];

   data_col116[1] <= data[49];
   data_col116[2] <= data_col116[1];
   data_col116[3] <= data_col116[2];
   data_col116[4] <= data_col116[3];
   data_col116[5] <= data_col116[4];
   data_col116[6] <= data_col116[5];
   data_col116[7] <= data_col116[6];
   data_col116[8] <= data_col116[7];
   data_col116[9] <= data_col116[8];
   data_col116[10] <= data_col116[9];
   data_col116[11] <= data_col116[10];
   data_col116[12] <= data_col116[11];
   data_col116[13] <= data_col116[12];
   data_col116[14] <= data_col116[13];
   data_col116[15] <= data_col116[14];
   data_col116[16] <= data_col116[15];
   data_col116[17] <= data_col116[16];
   data_col116[18] <= data_col116[17];
   data_col116[19] <= data_col116[18];
   data_col116[20] <= data_col116[19];
   data_col116[21] <= data_col116[20];
   data_col116[22] <= data_col116[21];
   data_col116[23] <= data_col116[22];
   data_col116[24] <= data_col116[23];
   data_col116[25] <= data_col116[24];
   data_col116[26] <= data_col116[25];
   data_col116[27] <= data_col116[26];
   data_col116[28] <= data_col116[27];
   data_col116[29] <= data_col116[28];
   data_col116[30] <= data_col116[29];
   data_col116[31] <= data_col116[30];
   data_col116[32] <= data_col116[31];
   data_col116[33] <= data_col116[32];
   data_col116[34] <= data_col116[33];
   data_col116[35] <= data_col116[34];
   data_col116[36] <= data_col116[35];
   data_col116[37] <= data_col116[36];
   data_col116[38] <= data_col116[37];
   data_col116[39] <= data_col116[38];
   data_col116[40] <= data_col116[39];
   data_col116[41] <= data_col116[40];
   data_col116[42] <= data_col116[41];
   data_col116[43] <= data_col116[42];
   data_col116[44] <= data_col116[43];
   data_col116[45] <= data_col116[44];
   data_col116[46] <= data_col116[45];
   data_col116[47] <= data_col116[46];
   data_col116[48] <= data_col116[47];
   data_col116[49] <= data_col116[48];
   data_col116[50] <= data_col116[49];
   data_col116[51] <= data_col116[50];
   data_col116[52] <= data_col116[51];
   data_col116[53] <= data_col116[52];
   data_col116[54] <= data_col116[53];
   data_col116[55] <= data_col116[54];
   data_col116[56] <= data_col116[55];
   data_col116[57] <= data_col116[56];
   data_col116[58] <= data_col116[57];
   data_col116[59] <= data_col116[58];
   data_col116[60] <= data_col116[59];
   data_col116[61] <= data_col116[60];
   data_col116[62] <= data_col116[61];
   data_col116[63] <= data_col116[62];
   data_col116[64] <= data_col116[63];
   data_col116[65] <= data_col116[64];
   data_col116[66] <= data_col116[65];
   data_col116[67] <= data_col116[66];
   data_col116[68] <= data_col116[67];
   data_col116[69] <= data_col116[68];
   data_col116[70] <= data_col116[69];
   data_col116[71] <= data_col116[70];
   data_col116[72] <= data_col116[71];
   data_col116[73] <= data_col116[72];
   data_col116[74] <= data_col116[73];
   data_col116[75] <= data_col116[74];
   data_col116[76] <= data_col116[75];
   data_col116[77] <= data_col116[76];
   data_col116[78] <= data_col116[77];
   data_col116[79] <= data_col116[78];
   data_col116[80] <= data_col116[79];
   data_col116[81] <= data_col116[80];
   data_col116[82] <= data_col116[81];
   data_col116[83] <= data_col116[82];
   data_col116[84] <= data_col116[83];
   data_col116[85] <= data_col116[84];
   data_col116[86] <= data_col116[85];
   data_col116[87] <= data_col116[86];
   data_col116[88] <= data_col116[87];
   data_col116[89] <= data_col116[88];
   data_col116[90] <= data_col116[89];
   data_col116[91] <= data_col116[90];
   data_col116[92] <= data_col116[91];
   data_col116[93] <= data_col116[92];
   data_col116[94] <= data_col116[93];
   data_col116[95] <= data_col116[94];
   data_col116[96] <= data_col116[95];
   data_col116[97] <= data_col116[96];
   data_col116[98] <= data_col116[97];
   data_col116[99] <= data_col116[98];
   data_col116[100] <= data_col116[99];
   data_col116[101] <= data_col116[100];
   data_col116[102] <= data_col116[101];
   data_col116[103] <= data_col116[102];
   data_col116[104] <= data_col116[103];
   data_col116[105] <= data_col116[104];
   data_col116[106] <= data_col116[105];
   data_col116[107] <= data_col116[106];
   data_col116[108] <= data_col116[107];
   data_col116[109] <= data_col116[108];
   data_col116[110] <= data_col116[109];
   data_col116[111] <= data_col116[110];
   data_col116[112] <= data_col116[111];
   data_col116[113] <= data_col116[112];
   data_col116[114] <= data_col116[113];
   data_col116[115] <= data_col116[114];
   data_col116[116] <= data_col116[115];

   data_col117[1] <= data[48];
   data_col117[2] <= data_col117[1];
   data_col117[3] <= data_col117[2];
   data_col117[4] <= data_col117[3];
   data_col117[5] <= data_col117[4];
   data_col117[6] <= data_col117[5];
   data_col117[7] <= data_col117[6];
   data_col117[8] <= data_col117[7];
   data_col117[9] <= data_col117[8];
   data_col117[10] <= data_col117[9];
   data_col117[11] <= data_col117[10];
   data_col117[12] <= data_col117[11];
   data_col117[13] <= data_col117[12];
   data_col117[14] <= data_col117[13];
   data_col117[15] <= data_col117[14];
   data_col117[16] <= data_col117[15];
   data_col117[17] <= data_col117[16];
   data_col117[18] <= data_col117[17];
   data_col117[19] <= data_col117[18];
   data_col117[20] <= data_col117[19];
   data_col117[21] <= data_col117[20];
   data_col117[22] <= data_col117[21];
   data_col117[23] <= data_col117[22];
   data_col117[24] <= data_col117[23];
   data_col117[25] <= data_col117[24];
   data_col117[26] <= data_col117[25];
   data_col117[27] <= data_col117[26];
   data_col117[28] <= data_col117[27];
   data_col117[29] <= data_col117[28];
   data_col117[30] <= data_col117[29];
   data_col117[31] <= data_col117[30];
   data_col117[32] <= data_col117[31];
   data_col117[33] <= data_col117[32];
   data_col117[34] <= data_col117[33];
   data_col117[35] <= data_col117[34];
   data_col117[36] <= data_col117[35];
   data_col117[37] <= data_col117[36];
   data_col117[38] <= data_col117[37];
   data_col117[39] <= data_col117[38];
   data_col117[40] <= data_col117[39];
   data_col117[41] <= data_col117[40];
   data_col117[42] <= data_col117[41];
   data_col117[43] <= data_col117[42];
   data_col117[44] <= data_col117[43];
   data_col117[45] <= data_col117[44];
   data_col117[46] <= data_col117[45];
   data_col117[47] <= data_col117[46];
   data_col117[48] <= data_col117[47];
   data_col117[49] <= data_col117[48];
   data_col117[50] <= data_col117[49];
   data_col117[51] <= data_col117[50];
   data_col117[52] <= data_col117[51];
   data_col117[53] <= data_col117[52];
   data_col117[54] <= data_col117[53];
   data_col117[55] <= data_col117[54];
   data_col117[56] <= data_col117[55];
   data_col117[57] <= data_col117[56];
   data_col117[58] <= data_col117[57];
   data_col117[59] <= data_col117[58];
   data_col117[60] <= data_col117[59];
   data_col117[61] <= data_col117[60];
   data_col117[62] <= data_col117[61];
   data_col117[63] <= data_col117[62];
   data_col117[64] <= data_col117[63];
   data_col117[65] <= data_col117[64];
   data_col117[66] <= data_col117[65];
   data_col117[67] <= data_col117[66];
   data_col117[68] <= data_col117[67];
   data_col117[69] <= data_col117[68];
   data_col117[70] <= data_col117[69];
   data_col117[71] <= data_col117[70];
   data_col117[72] <= data_col117[71];
   data_col117[73] <= data_col117[72];
   data_col117[74] <= data_col117[73];
   data_col117[75] <= data_col117[74];
   data_col117[76] <= data_col117[75];
   data_col117[77] <= data_col117[76];
   data_col117[78] <= data_col117[77];
   data_col117[79] <= data_col117[78];
   data_col117[80] <= data_col117[79];
   data_col117[81] <= data_col117[80];
   data_col117[82] <= data_col117[81];
   data_col117[83] <= data_col117[82];
   data_col117[84] <= data_col117[83];
   data_col117[85] <= data_col117[84];
   data_col117[86] <= data_col117[85];
   data_col117[87] <= data_col117[86];
   data_col117[88] <= data_col117[87];
   data_col117[89] <= data_col117[88];
   data_col117[90] <= data_col117[89];
   data_col117[91] <= data_col117[90];
   data_col117[92] <= data_col117[91];
   data_col117[93] <= data_col117[92];
   data_col117[94] <= data_col117[93];
   data_col117[95] <= data_col117[94];
   data_col117[96] <= data_col117[95];
   data_col117[97] <= data_col117[96];
   data_col117[98] <= data_col117[97];
   data_col117[99] <= data_col117[98];
   data_col117[100] <= data_col117[99];
   data_col117[101] <= data_col117[100];
   data_col117[102] <= data_col117[101];
   data_col117[103] <= data_col117[102];
   data_col117[104] <= data_col117[103];
   data_col117[105] <= data_col117[104];
   data_col117[106] <= data_col117[105];
   data_col117[107] <= data_col117[106];
   data_col117[108] <= data_col117[107];
   data_col117[109] <= data_col117[108];
   data_col117[110] <= data_col117[109];
   data_col117[111] <= data_col117[110];
   data_col117[112] <= data_col117[111];
   data_col117[113] <= data_col117[112];
   data_col117[114] <= data_col117[113];
   data_col117[115] <= data_col117[114];
   data_col117[116] <= data_col117[115];
   data_col117[117] <= data_col117[116];

   data_col118[1] <= data[47];
   data_col118[2] <= data_col118[1];
   data_col118[3] <= data_col118[2];
   data_col118[4] <= data_col118[3];
   data_col118[5] <= data_col118[4];
   data_col118[6] <= data_col118[5];
   data_col118[7] <= data_col118[6];
   data_col118[8] <= data_col118[7];
   data_col118[9] <= data_col118[8];
   data_col118[10] <= data_col118[9];
   data_col118[11] <= data_col118[10];
   data_col118[12] <= data_col118[11];
   data_col118[13] <= data_col118[12];
   data_col118[14] <= data_col118[13];
   data_col118[15] <= data_col118[14];
   data_col118[16] <= data_col118[15];
   data_col118[17] <= data_col118[16];
   data_col118[18] <= data_col118[17];
   data_col118[19] <= data_col118[18];
   data_col118[20] <= data_col118[19];
   data_col118[21] <= data_col118[20];
   data_col118[22] <= data_col118[21];
   data_col118[23] <= data_col118[22];
   data_col118[24] <= data_col118[23];
   data_col118[25] <= data_col118[24];
   data_col118[26] <= data_col118[25];
   data_col118[27] <= data_col118[26];
   data_col118[28] <= data_col118[27];
   data_col118[29] <= data_col118[28];
   data_col118[30] <= data_col118[29];
   data_col118[31] <= data_col118[30];
   data_col118[32] <= data_col118[31];
   data_col118[33] <= data_col118[32];
   data_col118[34] <= data_col118[33];
   data_col118[35] <= data_col118[34];
   data_col118[36] <= data_col118[35];
   data_col118[37] <= data_col118[36];
   data_col118[38] <= data_col118[37];
   data_col118[39] <= data_col118[38];
   data_col118[40] <= data_col118[39];
   data_col118[41] <= data_col118[40];
   data_col118[42] <= data_col118[41];
   data_col118[43] <= data_col118[42];
   data_col118[44] <= data_col118[43];
   data_col118[45] <= data_col118[44];
   data_col118[46] <= data_col118[45];
   data_col118[47] <= data_col118[46];
   data_col118[48] <= data_col118[47];
   data_col118[49] <= data_col118[48];
   data_col118[50] <= data_col118[49];
   data_col118[51] <= data_col118[50];
   data_col118[52] <= data_col118[51];
   data_col118[53] <= data_col118[52];
   data_col118[54] <= data_col118[53];
   data_col118[55] <= data_col118[54];
   data_col118[56] <= data_col118[55];
   data_col118[57] <= data_col118[56];
   data_col118[58] <= data_col118[57];
   data_col118[59] <= data_col118[58];
   data_col118[60] <= data_col118[59];
   data_col118[61] <= data_col118[60];
   data_col118[62] <= data_col118[61];
   data_col118[63] <= data_col118[62];
   data_col118[64] <= data_col118[63];
   data_col118[65] <= data_col118[64];
   data_col118[66] <= data_col118[65];
   data_col118[67] <= data_col118[66];
   data_col118[68] <= data_col118[67];
   data_col118[69] <= data_col118[68];
   data_col118[70] <= data_col118[69];
   data_col118[71] <= data_col118[70];
   data_col118[72] <= data_col118[71];
   data_col118[73] <= data_col118[72];
   data_col118[74] <= data_col118[73];
   data_col118[75] <= data_col118[74];
   data_col118[76] <= data_col118[75];
   data_col118[77] <= data_col118[76];
   data_col118[78] <= data_col118[77];
   data_col118[79] <= data_col118[78];
   data_col118[80] <= data_col118[79];
   data_col118[81] <= data_col118[80];
   data_col118[82] <= data_col118[81];
   data_col118[83] <= data_col118[82];
   data_col118[84] <= data_col118[83];
   data_col118[85] <= data_col118[84];
   data_col118[86] <= data_col118[85];
   data_col118[87] <= data_col118[86];
   data_col118[88] <= data_col118[87];
   data_col118[89] <= data_col118[88];
   data_col118[90] <= data_col118[89];
   data_col118[91] <= data_col118[90];
   data_col118[92] <= data_col118[91];
   data_col118[93] <= data_col118[92];
   data_col118[94] <= data_col118[93];
   data_col118[95] <= data_col118[94];
   data_col118[96] <= data_col118[95];
   data_col118[97] <= data_col118[96];
   data_col118[98] <= data_col118[97];
   data_col118[99] <= data_col118[98];
   data_col118[100] <= data_col118[99];
   data_col118[101] <= data_col118[100];
   data_col118[102] <= data_col118[101];
   data_col118[103] <= data_col118[102];
   data_col118[104] <= data_col118[103];
   data_col118[105] <= data_col118[104];
   data_col118[106] <= data_col118[105];
   data_col118[107] <= data_col118[106];
   data_col118[108] <= data_col118[107];
   data_col118[109] <= data_col118[108];
   data_col118[110] <= data_col118[109];
   data_col118[111] <= data_col118[110];
   data_col118[112] <= data_col118[111];
   data_col118[113] <= data_col118[112];
   data_col118[114] <= data_col118[113];
   data_col118[115] <= data_col118[114];
   data_col118[116] <= data_col118[115];
   data_col118[117] <= data_col118[116];
   data_col118[118] <= data_col118[117];

   data_col119[1] <= data[46];
   data_col119[2] <= data_col119[1];
   data_col119[3] <= data_col119[2];
   data_col119[4] <= data_col119[3];
   data_col119[5] <= data_col119[4];
   data_col119[6] <= data_col119[5];
   data_col119[7] <= data_col119[6];
   data_col119[8] <= data_col119[7];
   data_col119[9] <= data_col119[8];
   data_col119[10] <= data_col119[9];
   data_col119[11] <= data_col119[10];
   data_col119[12] <= data_col119[11];
   data_col119[13] <= data_col119[12];
   data_col119[14] <= data_col119[13];
   data_col119[15] <= data_col119[14];
   data_col119[16] <= data_col119[15];
   data_col119[17] <= data_col119[16];
   data_col119[18] <= data_col119[17];
   data_col119[19] <= data_col119[18];
   data_col119[20] <= data_col119[19];
   data_col119[21] <= data_col119[20];
   data_col119[22] <= data_col119[21];
   data_col119[23] <= data_col119[22];
   data_col119[24] <= data_col119[23];
   data_col119[25] <= data_col119[24];
   data_col119[26] <= data_col119[25];
   data_col119[27] <= data_col119[26];
   data_col119[28] <= data_col119[27];
   data_col119[29] <= data_col119[28];
   data_col119[30] <= data_col119[29];
   data_col119[31] <= data_col119[30];
   data_col119[32] <= data_col119[31];
   data_col119[33] <= data_col119[32];
   data_col119[34] <= data_col119[33];
   data_col119[35] <= data_col119[34];
   data_col119[36] <= data_col119[35];
   data_col119[37] <= data_col119[36];
   data_col119[38] <= data_col119[37];
   data_col119[39] <= data_col119[38];
   data_col119[40] <= data_col119[39];
   data_col119[41] <= data_col119[40];
   data_col119[42] <= data_col119[41];
   data_col119[43] <= data_col119[42];
   data_col119[44] <= data_col119[43];
   data_col119[45] <= data_col119[44];
   data_col119[46] <= data_col119[45];
   data_col119[47] <= data_col119[46];
   data_col119[48] <= data_col119[47];
   data_col119[49] <= data_col119[48];
   data_col119[50] <= data_col119[49];
   data_col119[51] <= data_col119[50];
   data_col119[52] <= data_col119[51];
   data_col119[53] <= data_col119[52];
   data_col119[54] <= data_col119[53];
   data_col119[55] <= data_col119[54];
   data_col119[56] <= data_col119[55];
   data_col119[57] <= data_col119[56];
   data_col119[58] <= data_col119[57];
   data_col119[59] <= data_col119[58];
   data_col119[60] <= data_col119[59];
   data_col119[61] <= data_col119[60];
   data_col119[62] <= data_col119[61];
   data_col119[63] <= data_col119[62];
   data_col119[64] <= data_col119[63];
   data_col119[65] <= data_col119[64];
   data_col119[66] <= data_col119[65];
   data_col119[67] <= data_col119[66];
   data_col119[68] <= data_col119[67];
   data_col119[69] <= data_col119[68];
   data_col119[70] <= data_col119[69];
   data_col119[71] <= data_col119[70];
   data_col119[72] <= data_col119[71];
   data_col119[73] <= data_col119[72];
   data_col119[74] <= data_col119[73];
   data_col119[75] <= data_col119[74];
   data_col119[76] <= data_col119[75];
   data_col119[77] <= data_col119[76];
   data_col119[78] <= data_col119[77];
   data_col119[79] <= data_col119[78];
   data_col119[80] <= data_col119[79];
   data_col119[81] <= data_col119[80];
   data_col119[82] <= data_col119[81];
   data_col119[83] <= data_col119[82];
   data_col119[84] <= data_col119[83];
   data_col119[85] <= data_col119[84];
   data_col119[86] <= data_col119[85];
   data_col119[87] <= data_col119[86];
   data_col119[88] <= data_col119[87];
   data_col119[89] <= data_col119[88];
   data_col119[90] <= data_col119[89];
   data_col119[91] <= data_col119[90];
   data_col119[92] <= data_col119[91];
   data_col119[93] <= data_col119[92];
   data_col119[94] <= data_col119[93];
   data_col119[95] <= data_col119[94];
   data_col119[96] <= data_col119[95];
   data_col119[97] <= data_col119[96];
   data_col119[98] <= data_col119[97];
   data_col119[99] <= data_col119[98];
   data_col119[100] <= data_col119[99];
   data_col119[101] <= data_col119[100];
   data_col119[102] <= data_col119[101];
   data_col119[103] <= data_col119[102];
   data_col119[104] <= data_col119[103];
   data_col119[105] <= data_col119[104];
   data_col119[106] <= data_col119[105];
   data_col119[107] <= data_col119[106];
   data_col119[108] <= data_col119[107];
   data_col119[109] <= data_col119[108];
   data_col119[110] <= data_col119[109];
   data_col119[111] <= data_col119[110];
   data_col119[112] <= data_col119[111];
   data_col119[113] <= data_col119[112];
   data_col119[114] <= data_col119[113];
   data_col119[115] <= data_col119[114];
   data_col119[116] <= data_col119[115];
   data_col119[117] <= data_col119[116];
   data_col119[118] <= data_col119[117];
   data_col119[119] <= data_col119[118];

   data_col120[1] <= data[45];
   data_col120[2] <= data_col120[1];
   data_col120[3] <= data_col120[2];
   data_col120[4] <= data_col120[3];
   data_col120[5] <= data_col120[4];
   data_col120[6] <= data_col120[5];
   data_col120[7] <= data_col120[6];
   data_col120[8] <= data_col120[7];
   data_col120[9] <= data_col120[8];
   data_col120[10] <= data_col120[9];
   data_col120[11] <= data_col120[10];
   data_col120[12] <= data_col120[11];
   data_col120[13] <= data_col120[12];
   data_col120[14] <= data_col120[13];
   data_col120[15] <= data_col120[14];
   data_col120[16] <= data_col120[15];
   data_col120[17] <= data_col120[16];
   data_col120[18] <= data_col120[17];
   data_col120[19] <= data_col120[18];
   data_col120[20] <= data_col120[19];
   data_col120[21] <= data_col120[20];
   data_col120[22] <= data_col120[21];
   data_col120[23] <= data_col120[22];
   data_col120[24] <= data_col120[23];
   data_col120[25] <= data_col120[24];
   data_col120[26] <= data_col120[25];
   data_col120[27] <= data_col120[26];
   data_col120[28] <= data_col120[27];
   data_col120[29] <= data_col120[28];
   data_col120[30] <= data_col120[29];
   data_col120[31] <= data_col120[30];
   data_col120[32] <= data_col120[31];
   data_col120[33] <= data_col120[32];
   data_col120[34] <= data_col120[33];
   data_col120[35] <= data_col120[34];
   data_col120[36] <= data_col120[35];
   data_col120[37] <= data_col120[36];
   data_col120[38] <= data_col120[37];
   data_col120[39] <= data_col120[38];
   data_col120[40] <= data_col120[39];
   data_col120[41] <= data_col120[40];
   data_col120[42] <= data_col120[41];
   data_col120[43] <= data_col120[42];
   data_col120[44] <= data_col120[43];
   data_col120[45] <= data_col120[44];
   data_col120[46] <= data_col120[45];
   data_col120[47] <= data_col120[46];
   data_col120[48] <= data_col120[47];
   data_col120[49] <= data_col120[48];
   data_col120[50] <= data_col120[49];
   data_col120[51] <= data_col120[50];
   data_col120[52] <= data_col120[51];
   data_col120[53] <= data_col120[52];
   data_col120[54] <= data_col120[53];
   data_col120[55] <= data_col120[54];
   data_col120[56] <= data_col120[55];
   data_col120[57] <= data_col120[56];
   data_col120[58] <= data_col120[57];
   data_col120[59] <= data_col120[58];
   data_col120[60] <= data_col120[59];
   data_col120[61] <= data_col120[60];
   data_col120[62] <= data_col120[61];
   data_col120[63] <= data_col120[62];
   data_col120[64] <= data_col120[63];
   data_col120[65] <= data_col120[64];
   data_col120[66] <= data_col120[65];
   data_col120[67] <= data_col120[66];
   data_col120[68] <= data_col120[67];
   data_col120[69] <= data_col120[68];
   data_col120[70] <= data_col120[69];
   data_col120[71] <= data_col120[70];
   data_col120[72] <= data_col120[71];
   data_col120[73] <= data_col120[72];
   data_col120[74] <= data_col120[73];
   data_col120[75] <= data_col120[74];
   data_col120[76] <= data_col120[75];
   data_col120[77] <= data_col120[76];
   data_col120[78] <= data_col120[77];
   data_col120[79] <= data_col120[78];
   data_col120[80] <= data_col120[79];
   data_col120[81] <= data_col120[80];
   data_col120[82] <= data_col120[81];
   data_col120[83] <= data_col120[82];
   data_col120[84] <= data_col120[83];
   data_col120[85] <= data_col120[84];
   data_col120[86] <= data_col120[85];
   data_col120[87] <= data_col120[86];
   data_col120[88] <= data_col120[87];
   data_col120[89] <= data_col120[88];
   data_col120[90] <= data_col120[89];
   data_col120[91] <= data_col120[90];
   data_col120[92] <= data_col120[91];
   data_col120[93] <= data_col120[92];
   data_col120[94] <= data_col120[93];
   data_col120[95] <= data_col120[94];
   data_col120[96] <= data_col120[95];
   data_col120[97] <= data_col120[96];
   data_col120[98] <= data_col120[97];
   data_col120[99] <= data_col120[98];
   data_col120[100] <= data_col120[99];
   data_col120[101] <= data_col120[100];
   data_col120[102] <= data_col120[101];
   data_col120[103] <= data_col120[102];
   data_col120[104] <= data_col120[103];
   data_col120[105] <= data_col120[104];
   data_col120[106] <= data_col120[105];
   data_col120[107] <= data_col120[106];
   data_col120[108] <= data_col120[107];
   data_col120[109] <= data_col120[108];
   data_col120[110] <= data_col120[109];
   data_col120[111] <= data_col120[110];
   data_col120[112] <= data_col120[111];
   data_col120[113] <= data_col120[112];
   data_col120[114] <= data_col120[113];
   data_col120[115] <= data_col120[114];
   data_col120[116] <= data_col120[115];
   data_col120[117] <= data_col120[116];
   data_col120[118] <= data_col120[117];
   data_col120[119] <= data_col120[118];
   data_col120[120] <= data_col120[119];

   data_col121[1] <= data[44];
   data_col121[2] <= data_col121[1];
   data_col121[3] <= data_col121[2];
   data_col121[4] <= data_col121[3];
   data_col121[5] <= data_col121[4];
   data_col121[6] <= data_col121[5];
   data_col121[7] <= data_col121[6];
   data_col121[8] <= data_col121[7];
   data_col121[9] <= data_col121[8];
   data_col121[10] <= data_col121[9];
   data_col121[11] <= data_col121[10];
   data_col121[12] <= data_col121[11];
   data_col121[13] <= data_col121[12];
   data_col121[14] <= data_col121[13];
   data_col121[15] <= data_col121[14];
   data_col121[16] <= data_col121[15];
   data_col121[17] <= data_col121[16];
   data_col121[18] <= data_col121[17];
   data_col121[19] <= data_col121[18];
   data_col121[20] <= data_col121[19];
   data_col121[21] <= data_col121[20];
   data_col121[22] <= data_col121[21];
   data_col121[23] <= data_col121[22];
   data_col121[24] <= data_col121[23];
   data_col121[25] <= data_col121[24];
   data_col121[26] <= data_col121[25];
   data_col121[27] <= data_col121[26];
   data_col121[28] <= data_col121[27];
   data_col121[29] <= data_col121[28];
   data_col121[30] <= data_col121[29];
   data_col121[31] <= data_col121[30];
   data_col121[32] <= data_col121[31];
   data_col121[33] <= data_col121[32];
   data_col121[34] <= data_col121[33];
   data_col121[35] <= data_col121[34];
   data_col121[36] <= data_col121[35];
   data_col121[37] <= data_col121[36];
   data_col121[38] <= data_col121[37];
   data_col121[39] <= data_col121[38];
   data_col121[40] <= data_col121[39];
   data_col121[41] <= data_col121[40];
   data_col121[42] <= data_col121[41];
   data_col121[43] <= data_col121[42];
   data_col121[44] <= data_col121[43];
   data_col121[45] <= data_col121[44];
   data_col121[46] <= data_col121[45];
   data_col121[47] <= data_col121[46];
   data_col121[48] <= data_col121[47];
   data_col121[49] <= data_col121[48];
   data_col121[50] <= data_col121[49];
   data_col121[51] <= data_col121[50];
   data_col121[52] <= data_col121[51];
   data_col121[53] <= data_col121[52];
   data_col121[54] <= data_col121[53];
   data_col121[55] <= data_col121[54];
   data_col121[56] <= data_col121[55];
   data_col121[57] <= data_col121[56];
   data_col121[58] <= data_col121[57];
   data_col121[59] <= data_col121[58];
   data_col121[60] <= data_col121[59];
   data_col121[61] <= data_col121[60];
   data_col121[62] <= data_col121[61];
   data_col121[63] <= data_col121[62];
   data_col121[64] <= data_col121[63];
   data_col121[65] <= data_col121[64];
   data_col121[66] <= data_col121[65];
   data_col121[67] <= data_col121[66];
   data_col121[68] <= data_col121[67];
   data_col121[69] <= data_col121[68];
   data_col121[70] <= data_col121[69];
   data_col121[71] <= data_col121[70];
   data_col121[72] <= data_col121[71];
   data_col121[73] <= data_col121[72];
   data_col121[74] <= data_col121[73];
   data_col121[75] <= data_col121[74];
   data_col121[76] <= data_col121[75];
   data_col121[77] <= data_col121[76];
   data_col121[78] <= data_col121[77];
   data_col121[79] <= data_col121[78];
   data_col121[80] <= data_col121[79];
   data_col121[81] <= data_col121[80];
   data_col121[82] <= data_col121[81];
   data_col121[83] <= data_col121[82];
   data_col121[84] <= data_col121[83];
   data_col121[85] <= data_col121[84];
   data_col121[86] <= data_col121[85];
   data_col121[87] <= data_col121[86];
   data_col121[88] <= data_col121[87];
   data_col121[89] <= data_col121[88];
   data_col121[90] <= data_col121[89];
   data_col121[91] <= data_col121[90];
   data_col121[92] <= data_col121[91];
   data_col121[93] <= data_col121[92];
   data_col121[94] <= data_col121[93];
   data_col121[95] <= data_col121[94];
   data_col121[96] <= data_col121[95];
   data_col121[97] <= data_col121[96];
   data_col121[98] <= data_col121[97];
   data_col121[99] <= data_col121[98];
   data_col121[100] <= data_col121[99];
   data_col121[101] <= data_col121[100];
   data_col121[102] <= data_col121[101];
   data_col121[103] <= data_col121[102];
   data_col121[104] <= data_col121[103];
   data_col121[105] <= data_col121[104];
   data_col121[106] <= data_col121[105];
   data_col121[107] <= data_col121[106];
   data_col121[108] <= data_col121[107];
   data_col121[109] <= data_col121[108];
   data_col121[110] <= data_col121[109];
   data_col121[111] <= data_col121[110];
   data_col121[112] <= data_col121[111];
   data_col121[113] <= data_col121[112];
   data_col121[114] <= data_col121[113];
   data_col121[115] <= data_col121[114];
   data_col121[116] <= data_col121[115];
   data_col121[117] <= data_col121[116];
   data_col121[118] <= data_col121[117];
   data_col121[119] <= data_col121[118];
   data_col121[120] <= data_col121[119];
   data_col121[121] <= data_col121[120];

   data_col122[1] <= data[43];
   data_col122[2] <= data_col122[1];
   data_col122[3] <= data_col122[2];
   data_col122[4] <= data_col122[3];
   data_col122[5] <= data_col122[4];
   data_col122[6] <= data_col122[5];
   data_col122[7] <= data_col122[6];
   data_col122[8] <= data_col122[7];
   data_col122[9] <= data_col122[8];
   data_col122[10] <= data_col122[9];
   data_col122[11] <= data_col122[10];
   data_col122[12] <= data_col122[11];
   data_col122[13] <= data_col122[12];
   data_col122[14] <= data_col122[13];
   data_col122[15] <= data_col122[14];
   data_col122[16] <= data_col122[15];
   data_col122[17] <= data_col122[16];
   data_col122[18] <= data_col122[17];
   data_col122[19] <= data_col122[18];
   data_col122[20] <= data_col122[19];
   data_col122[21] <= data_col122[20];
   data_col122[22] <= data_col122[21];
   data_col122[23] <= data_col122[22];
   data_col122[24] <= data_col122[23];
   data_col122[25] <= data_col122[24];
   data_col122[26] <= data_col122[25];
   data_col122[27] <= data_col122[26];
   data_col122[28] <= data_col122[27];
   data_col122[29] <= data_col122[28];
   data_col122[30] <= data_col122[29];
   data_col122[31] <= data_col122[30];
   data_col122[32] <= data_col122[31];
   data_col122[33] <= data_col122[32];
   data_col122[34] <= data_col122[33];
   data_col122[35] <= data_col122[34];
   data_col122[36] <= data_col122[35];
   data_col122[37] <= data_col122[36];
   data_col122[38] <= data_col122[37];
   data_col122[39] <= data_col122[38];
   data_col122[40] <= data_col122[39];
   data_col122[41] <= data_col122[40];
   data_col122[42] <= data_col122[41];
   data_col122[43] <= data_col122[42];
   data_col122[44] <= data_col122[43];
   data_col122[45] <= data_col122[44];
   data_col122[46] <= data_col122[45];
   data_col122[47] <= data_col122[46];
   data_col122[48] <= data_col122[47];
   data_col122[49] <= data_col122[48];
   data_col122[50] <= data_col122[49];
   data_col122[51] <= data_col122[50];
   data_col122[52] <= data_col122[51];
   data_col122[53] <= data_col122[52];
   data_col122[54] <= data_col122[53];
   data_col122[55] <= data_col122[54];
   data_col122[56] <= data_col122[55];
   data_col122[57] <= data_col122[56];
   data_col122[58] <= data_col122[57];
   data_col122[59] <= data_col122[58];
   data_col122[60] <= data_col122[59];
   data_col122[61] <= data_col122[60];
   data_col122[62] <= data_col122[61];
   data_col122[63] <= data_col122[62];
   data_col122[64] <= data_col122[63];
   data_col122[65] <= data_col122[64];
   data_col122[66] <= data_col122[65];
   data_col122[67] <= data_col122[66];
   data_col122[68] <= data_col122[67];
   data_col122[69] <= data_col122[68];
   data_col122[70] <= data_col122[69];
   data_col122[71] <= data_col122[70];
   data_col122[72] <= data_col122[71];
   data_col122[73] <= data_col122[72];
   data_col122[74] <= data_col122[73];
   data_col122[75] <= data_col122[74];
   data_col122[76] <= data_col122[75];
   data_col122[77] <= data_col122[76];
   data_col122[78] <= data_col122[77];
   data_col122[79] <= data_col122[78];
   data_col122[80] <= data_col122[79];
   data_col122[81] <= data_col122[80];
   data_col122[82] <= data_col122[81];
   data_col122[83] <= data_col122[82];
   data_col122[84] <= data_col122[83];
   data_col122[85] <= data_col122[84];
   data_col122[86] <= data_col122[85];
   data_col122[87] <= data_col122[86];
   data_col122[88] <= data_col122[87];
   data_col122[89] <= data_col122[88];
   data_col122[90] <= data_col122[89];
   data_col122[91] <= data_col122[90];
   data_col122[92] <= data_col122[91];
   data_col122[93] <= data_col122[92];
   data_col122[94] <= data_col122[93];
   data_col122[95] <= data_col122[94];
   data_col122[96] <= data_col122[95];
   data_col122[97] <= data_col122[96];
   data_col122[98] <= data_col122[97];
   data_col122[99] <= data_col122[98];
   data_col122[100] <= data_col122[99];
   data_col122[101] <= data_col122[100];
   data_col122[102] <= data_col122[101];
   data_col122[103] <= data_col122[102];
   data_col122[104] <= data_col122[103];
   data_col122[105] <= data_col122[104];
   data_col122[106] <= data_col122[105];
   data_col122[107] <= data_col122[106];
   data_col122[108] <= data_col122[107];
   data_col122[109] <= data_col122[108];
   data_col122[110] <= data_col122[109];
   data_col122[111] <= data_col122[110];
   data_col122[112] <= data_col122[111];
   data_col122[113] <= data_col122[112];
   data_col122[114] <= data_col122[113];
   data_col122[115] <= data_col122[114];
   data_col122[116] <= data_col122[115];
   data_col122[117] <= data_col122[116];
   data_col122[118] <= data_col122[117];
   data_col122[119] <= data_col122[118];
   data_col122[120] <= data_col122[119];
   data_col122[121] <= data_col122[120];
   data_col122[122] <= data_col122[121];

   data_col123[1] <= data[42];
   data_col123[2] <= data_col123[1];
   data_col123[3] <= data_col123[2];
   data_col123[4] <= data_col123[3];
   data_col123[5] <= data_col123[4];
   data_col123[6] <= data_col123[5];
   data_col123[7] <= data_col123[6];
   data_col123[8] <= data_col123[7];
   data_col123[9] <= data_col123[8];
   data_col123[10] <= data_col123[9];
   data_col123[11] <= data_col123[10];
   data_col123[12] <= data_col123[11];
   data_col123[13] <= data_col123[12];
   data_col123[14] <= data_col123[13];
   data_col123[15] <= data_col123[14];
   data_col123[16] <= data_col123[15];
   data_col123[17] <= data_col123[16];
   data_col123[18] <= data_col123[17];
   data_col123[19] <= data_col123[18];
   data_col123[20] <= data_col123[19];
   data_col123[21] <= data_col123[20];
   data_col123[22] <= data_col123[21];
   data_col123[23] <= data_col123[22];
   data_col123[24] <= data_col123[23];
   data_col123[25] <= data_col123[24];
   data_col123[26] <= data_col123[25];
   data_col123[27] <= data_col123[26];
   data_col123[28] <= data_col123[27];
   data_col123[29] <= data_col123[28];
   data_col123[30] <= data_col123[29];
   data_col123[31] <= data_col123[30];
   data_col123[32] <= data_col123[31];
   data_col123[33] <= data_col123[32];
   data_col123[34] <= data_col123[33];
   data_col123[35] <= data_col123[34];
   data_col123[36] <= data_col123[35];
   data_col123[37] <= data_col123[36];
   data_col123[38] <= data_col123[37];
   data_col123[39] <= data_col123[38];
   data_col123[40] <= data_col123[39];
   data_col123[41] <= data_col123[40];
   data_col123[42] <= data_col123[41];
   data_col123[43] <= data_col123[42];
   data_col123[44] <= data_col123[43];
   data_col123[45] <= data_col123[44];
   data_col123[46] <= data_col123[45];
   data_col123[47] <= data_col123[46];
   data_col123[48] <= data_col123[47];
   data_col123[49] <= data_col123[48];
   data_col123[50] <= data_col123[49];
   data_col123[51] <= data_col123[50];
   data_col123[52] <= data_col123[51];
   data_col123[53] <= data_col123[52];
   data_col123[54] <= data_col123[53];
   data_col123[55] <= data_col123[54];
   data_col123[56] <= data_col123[55];
   data_col123[57] <= data_col123[56];
   data_col123[58] <= data_col123[57];
   data_col123[59] <= data_col123[58];
   data_col123[60] <= data_col123[59];
   data_col123[61] <= data_col123[60];
   data_col123[62] <= data_col123[61];
   data_col123[63] <= data_col123[62];
   data_col123[64] <= data_col123[63];
   data_col123[65] <= data_col123[64];
   data_col123[66] <= data_col123[65];
   data_col123[67] <= data_col123[66];
   data_col123[68] <= data_col123[67];
   data_col123[69] <= data_col123[68];
   data_col123[70] <= data_col123[69];
   data_col123[71] <= data_col123[70];
   data_col123[72] <= data_col123[71];
   data_col123[73] <= data_col123[72];
   data_col123[74] <= data_col123[73];
   data_col123[75] <= data_col123[74];
   data_col123[76] <= data_col123[75];
   data_col123[77] <= data_col123[76];
   data_col123[78] <= data_col123[77];
   data_col123[79] <= data_col123[78];
   data_col123[80] <= data_col123[79];
   data_col123[81] <= data_col123[80];
   data_col123[82] <= data_col123[81];
   data_col123[83] <= data_col123[82];
   data_col123[84] <= data_col123[83];
   data_col123[85] <= data_col123[84];
   data_col123[86] <= data_col123[85];
   data_col123[87] <= data_col123[86];
   data_col123[88] <= data_col123[87];
   data_col123[89] <= data_col123[88];
   data_col123[90] <= data_col123[89];
   data_col123[91] <= data_col123[90];
   data_col123[92] <= data_col123[91];
   data_col123[93] <= data_col123[92];
   data_col123[94] <= data_col123[93];
   data_col123[95] <= data_col123[94];
   data_col123[96] <= data_col123[95];
   data_col123[97] <= data_col123[96];
   data_col123[98] <= data_col123[97];
   data_col123[99] <= data_col123[98];
   data_col123[100] <= data_col123[99];
   data_col123[101] <= data_col123[100];
   data_col123[102] <= data_col123[101];
   data_col123[103] <= data_col123[102];
   data_col123[104] <= data_col123[103];
   data_col123[105] <= data_col123[104];
   data_col123[106] <= data_col123[105];
   data_col123[107] <= data_col123[106];
   data_col123[108] <= data_col123[107];
   data_col123[109] <= data_col123[108];
   data_col123[110] <= data_col123[109];
   data_col123[111] <= data_col123[110];
   data_col123[112] <= data_col123[111];
   data_col123[113] <= data_col123[112];
   data_col123[114] <= data_col123[113];
   data_col123[115] <= data_col123[114];
   data_col123[116] <= data_col123[115];
   data_col123[117] <= data_col123[116];
   data_col123[118] <= data_col123[117];
   data_col123[119] <= data_col123[118];
   data_col123[120] <= data_col123[119];
   data_col123[121] <= data_col123[120];
   data_col123[122] <= data_col123[121];
   data_col123[123] <= data_col123[122];

   data_col124[1] <= data[41];
   data_col124[2] <= data_col124[1];
   data_col124[3] <= data_col124[2];
   data_col124[4] <= data_col124[3];
   data_col124[5] <= data_col124[4];
   data_col124[6] <= data_col124[5];
   data_col124[7] <= data_col124[6];
   data_col124[8] <= data_col124[7];
   data_col124[9] <= data_col124[8];
   data_col124[10] <= data_col124[9];
   data_col124[11] <= data_col124[10];
   data_col124[12] <= data_col124[11];
   data_col124[13] <= data_col124[12];
   data_col124[14] <= data_col124[13];
   data_col124[15] <= data_col124[14];
   data_col124[16] <= data_col124[15];
   data_col124[17] <= data_col124[16];
   data_col124[18] <= data_col124[17];
   data_col124[19] <= data_col124[18];
   data_col124[20] <= data_col124[19];
   data_col124[21] <= data_col124[20];
   data_col124[22] <= data_col124[21];
   data_col124[23] <= data_col124[22];
   data_col124[24] <= data_col124[23];
   data_col124[25] <= data_col124[24];
   data_col124[26] <= data_col124[25];
   data_col124[27] <= data_col124[26];
   data_col124[28] <= data_col124[27];
   data_col124[29] <= data_col124[28];
   data_col124[30] <= data_col124[29];
   data_col124[31] <= data_col124[30];
   data_col124[32] <= data_col124[31];
   data_col124[33] <= data_col124[32];
   data_col124[34] <= data_col124[33];
   data_col124[35] <= data_col124[34];
   data_col124[36] <= data_col124[35];
   data_col124[37] <= data_col124[36];
   data_col124[38] <= data_col124[37];
   data_col124[39] <= data_col124[38];
   data_col124[40] <= data_col124[39];
   data_col124[41] <= data_col124[40];
   data_col124[42] <= data_col124[41];
   data_col124[43] <= data_col124[42];
   data_col124[44] <= data_col124[43];
   data_col124[45] <= data_col124[44];
   data_col124[46] <= data_col124[45];
   data_col124[47] <= data_col124[46];
   data_col124[48] <= data_col124[47];
   data_col124[49] <= data_col124[48];
   data_col124[50] <= data_col124[49];
   data_col124[51] <= data_col124[50];
   data_col124[52] <= data_col124[51];
   data_col124[53] <= data_col124[52];
   data_col124[54] <= data_col124[53];
   data_col124[55] <= data_col124[54];
   data_col124[56] <= data_col124[55];
   data_col124[57] <= data_col124[56];
   data_col124[58] <= data_col124[57];
   data_col124[59] <= data_col124[58];
   data_col124[60] <= data_col124[59];
   data_col124[61] <= data_col124[60];
   data_col124[62] <= data_col124[61];
   data_col124[63] <= data_col124[62];
   data_col124[64] <= data_col124[63];
   data_col124[65] <= data_col124[64];
   data_col124[66] <= data_col124[65];
   data_col124[67] <= data_col124[66];
   data_col124[68] <= data_col124[67];
   data_col124[69] <= data_col124[68];
   data_col124[70] <= data_col124[69];
   data_col124[71] <= data_col124[70];
   data_col124[72] <= data_col124[71];
   data_col124[73] <= data_col124[72];
   data_col124[74] <= data_col124[73];
   data_col124[75] <= data_col124[74];
   data_col124[76] <= data_col124[75];
   data_col124[77] <= data_col124[76];
   data_col124[78] <= data_col124[77];
   data_col124[79] <= data_col124[78];
   data_col124[80] <= data_col124[79];
   data_col124[81] <= data_col124[80];
   data_col124[82] <= data_col124[81];
   data_col124[83] <= data_col124[82];
   data_col124[84] <= data_col124[83];
   data_col124[85] <= data_col124[84];
   data_col124[86] <= data_col124[85];
   data_col124[87] <= data_col124[86];
   data_col124[88] <= data_col124[87];
   data_col124[89] <= data_col124[88];
   data_col124[90] <= data_col124[89];
   data_col124[91] <= data_col124[90];
   data_col124[92] <= data_col124[91];
   data_col124[93] <= data_col124[92];
   data_col124[94] <= data_col124[93];
   data_col124[95] <= data_col124[94];
   data_col124[96] <= data_col124[95];
   data_col124[97] <= data_col124[96];
   data_col124[98] <= data_col124[97];
   data_col124[99] <= data_col124[98];
   data_col124[100] <= data_col124[99];
   data_col124[101] <= data_col124[100];
   data_col124[102] <= data_col124[101];
   data_col124[103] <= data_col124[102];
   data_col124[104] <= data_col124[103];
   data_col124[105] <= data_col124[104];
   data_col124[106] <= data_col124[105];
   data_col124[107] <= data_col124[106];
   data_col124[108] <= data_col124[107];
   data_col124[109] <= data_col124[108];
   data_col124[110] <= data_col124[109];
   data_col124[111] <= data_col124[110];
   data_col124[112] <= data_col124[111];
   data_col124[113] <= data_col124[112];
   data_col124[114] <= data_col124[113];
   data_col124[115] <= data_col124[114];
   data_col124[116] <= data_col124[115];
   data_col124[117] <= data_col124[116];
   data_col124[118] <= data_col124[117];
   data_col124[119] <= data_col124[118];
   data_col124[120] <= data_col124[119];
   data_col124[121] <= data_col124[120];
   data_col124[122] <= data_col124[121];
   data_col124[123] <= data_col124[122];
   data_col124[124] <= data_col124[123];

   data_col125[1] <= data[40];
   data_col125[2] <= data_col125[1];
   data_col125[3] <= data_col125[2];
   data_col125[4] <= data_col125[3];
   data_col125[5] <= data_col125[4];
   data_col125[6] <= data_col125[5];
   data_col125[7] <= data_col125[6];
   data_col125[8] <= data_col125[7];
   data_col125[9] <= data_col125[8];
   data_col125[10] <= data_col125[9];
   data_col125[11] <= data_col125[10];
   data_col125[12] <= data_col125[11];
   data_col125[13] <= data_col125[12];
   data_col125[14] <= data_col125[13];
   data_col125[15] <= data_col125[14];
   data_col125[16] <= data_col125[15];
   data_col125[17] <= data_col125[16];
   data_col125[18] <= data_col125[17];
   data_col125[19] <= data_col125[18];
   data_col125[20] <= data_col125[19];
   data_col125[21] <= data_col125[20];
   data_col125[22] <= data_col125[21];
   data_col125[23] <= data_col125[22];
   data_col125[24] <= data_col125[23];
   data_col125[25] <= data_col125[24];
   data_col125[26] <= data_col125[25];
   data_col125[27] <= data_col125[26];
   data_col125[28] <= data_col125[27];
   data_col125[29] <= data_col125[28];
   data_col125[30] <= data_col125[29];
   data_col125[31] <= data_col125[30];
   data_col125[32] <= data_col125[31];
   data_col125[33] <= data_col125[32];
   data_col125[34] <= data_col125[33];
   data_col125[35] <= data_col125[34];
   data_col125[36] <= data_col125[35];
   data_col125[37] <= data_col125[36];
   data_col125[38] <= data_col125[37];
   data_col125[39] <= data_col125[38];
   data_col125[40] <= data_col125[39];
   data_col125[41] <= data_col125[40];
   data_col125[42] <= data_col125[41];
   data_col125[43] <= data_col125[42];
   data_col125[44] <= data_col125[43];
   data_col125[45] <= data_col125[44];
   data_col125[46] <= data_col125[45];
   data_col125[47] <= data_col125[46];
   data_col125[48] <= data_col125[47];
   data_col125[49] <= data_col125[48];
   data_col125[50] <= data_col125[49];
   data_col125[51] <= data_col125[50];
   data_col125[52] <= data_col125[51];
   data_col125[53] <= data_col125[52];
   data_col125[54] <= data_col125[53];
   data_col125[55] <= data_col125[54];
   data_col125[56] <= data_col125[55];
   data_col125[57] <= data_col125[56];
   data_col125[58] <= data_col125[57];
   data_col125[59] <= data_col125[58];
   data_col125[60] <= data_col125[59];
   data_col125[61] <= data_col125[60];
   data_col125[62] <= data_col125[61];
   data_col125[63] <= data_col125[62];
   data_col125[64] <= data_col125[63];
   data_col125[65] <= data_col125[64];
   data_col125[66] <= data_col125[65];
   data_col125[67] <= data_col125[66];
   data_col125[68] <= data_col125[67];
   data_col125[69] <= data_col125[68];
   data_col125[70] <= data_col125[69];
   data_col125[71] <= data_col125[70];
   data_col125[72] <= data_col125[71];
   data_col125[73] <= data_col125[72];
   data_col125[74] <= data_col125[73];
   data_col125[75] <= data_col125[74];
   data_col125[76] <= data_col125[75];
   data_col125[77] <= data_col125[76];
   data_col125[78] <= data_col125[77];
   data_col125[79] <= data_col125[78];
   data_col125[80] <= data_col125[79];
   data_col125[81] <= data_col125[80];
   data_col125[82] <= data_col125[81];
   data_col125[83] <= data_col125[82];
   data_col125[84] <= data_col125[83];
   data_col125[85] <= data_col125[84];
   data_col125[86] <= data_col125[85];
   data_col125[87] <= data_col125[86];
   data_col125[88] <= data_col125[87];
   data_col125[89] <= data_col125[88];
   data_col125[90] <= data_col125[89];
   data_col125[91] <= data_col125[90];
   data_col125[92] <= data_col125[91];
   data_col125[93] <= data_col125[92];
   data_col125[94] <= data_col125[93];
   data_col125[95] <= data_col125[94];
   data_col125[96] <= data_col125[95];
   data_col125[97] <= data_col125[96];
   data_col125[98] <= data_col125[97];
   data_col125[99] <= data_col125[98];
   data_col125[100] <= data_col125[99];
   data_col125[101] <= data_col125[100];
   data_col125[102] <= data_col125[101];
   data_col125[103] <= data_col125[102];
   data_col125[104] <= data_col125[103];
   data_col125[105] <= data_col125[104];
   data_col125[106] <= data_col125[105];
   data_col125[107] <= data_col125[106];
   data_col125[108] <= data_col125[107];
   data_col125[109] <= data_col125[108];
   data_col125[110] <= data_col125[109];
   data_col125[111] <= data_col125[110];
   data_col125[112] <= data_col125[111];
   data_col125[113] <= data_col125[112];
   data_col125[114] <= data_col125[113];
   data_col125[115] <= data_col125[114];
   data_col125[116] <= data_col125[115];
   data_col125[117] <= data_col125[116];
   data_col125[118] <= data_col125[117];
   data_col125[119] <= data_col125[118];
   data_col125[120] <= data_col125[119];
   data_col125[121] <= data_col125[120];
   data_col125[122] <= data_col125[121];
   data_col125[123] <= data_col125[122];
   data_col125[124] <= data_col125[123];
   data_col125[125] <= data_col125[124];

   data_col126[1] <= data[39];
   data_col126[2] <= data_col126[1];
   data_col126[3] <= data_col126[2];
   data_col126[4] <= data_col126[3];
   data_col126[5] <= data_col126[4];
   data_col126[6] <= data_col126[5];
   data_col126[7] <= data_col126[6];
   data_col126[8] <= data_col126[7];
   data_col126[9] <= data_col126[8];
   data_col126[10] <= data_col126[9];
   data_col126[11] <= data_col126[10];
   data_col126[12] <= data_col126[11];
   data_col126[13] <= data_col126[12];
   data_col126[14] <= data_col126[13];
   data_col126[15] <= data_col126[14];
   data_col126[16] <= data_col126[15];
   data_col126[17] <= data_col126[16];
   data_col126[18] <= data_col126[17];
   data_col126[19] <= data_col126[18];
   data_col126[20] <= data_col126[19];
   data_col126[21] <= data_col126[20];
   data_col126[22] <= data_col126[21];
   data_col126[23] <= data_col126[22];
   data_col126[24] <= data_col126[23];
   data_col126[25] <= data_col126[24];
   data_col126[26] <= data_col126[25];
   data_col126[27] <= data_col126[26];
   data_col126[28] <= data_col126[27];
   data_col126[29] <= data_col126[28];
   data_col126[30] <= data_col126[29];
   data_col126[31] <= data_col126[30];
   data_col126[32] <= data_col126[31];
   data_col126[33] <= data_col126[32];
   data_col126[34] <= data_col126[33];
   data_col126[35] <= data_col126[34];
   data_col126[36] <= data_col126[35];
   data_col126[37] <= data_col126[36];
   data_col126[38] <= data_col126[37];
   data_col126[39] <= data_col126[38];
   data_col126[40] <= data_col126[39];
   data_col126[41] <= data_col126[40];
   data_col126[42] <= data_col126[41];
   data_col126[43] <= data_col126[42];
   data_col126[44] <= data_col126[43];
   data_col126[45] <= data_col126[44];
   data_col126[46] <= data_col126[45];
   data_col126[47] <= data_col126[46];
   data_col126[48] <= data_col126[47];
   data_col126[49] <= data_col126[48];
   data_col126[50] <= data_col126[49];
   data_col126[51] <= data_col126[50];
   data_col126[52] <= data_col126[51];
   data_col126[53] <= data_col126[52];
   data_col126[54] <= data_col126[53];
   data_col126[55] <= data_col126[54];
   data_col126[56] <= data_col126[55];
   data_col126[57] <= data_col126[56];
   data_col126[58] <= data_col126[57];
   data_col126[59] <= data_col126[58];
   data_col126[60] <= data_col126[59];
   data_col126[61] <= data_col126[60];
   data_col126[62] <= data_col126[61];
   data_col126[63] <= data_col126[62];
   data_col126[64] <= data_col126[63];
   data_col126[65] <= data_col126[64];
   data_col126[66] <= data_col126[65];
   data_col126[67] <= data_col126[66];
   data_col126[68] <= data_col126[67];
   data_col126[69] <= data_col126[68];
   data_col126[70] <= data_col126[69];
   data_col126[71] <= data_col126[70];
   data_col126[72] <= data_col126[71];
   data_col126[73] <= data_col126[72];
   data_col126[74] <= data_col126[73];
   data_col126[75] <= data_col126[74];
   data_col126[76] <= data_col126[75];
   data_col126[77] <= data_col126[76];
   data_col126[78] <= data_col126[77];
   data_col126[79] <= data_col126[78];
   data_col126[80] <= data_col126[79];
   data_col126[81] <= data_col126[80];
   data_col126[82] <= data_col126[81];
   data_col126[83] <= data_col126[82];
   data_col126[84] <= data_col126[83];
   data_col126[85] <= data_col126[84];
   data_col126[86] <= data_col126[85];
   data_col126[87] <= data_col126[86];
   data_col126[88] <= data_col126[87];
   data_col126[89] <= data_col126[88];
   data_col126[90] <= data_col126[89];
   data_col126[91] <= data_col126[90];
   data_col126[92] <= data_col126[91];
   data_col126[93] <= data_col126[92];
   data_col126[94] <= data_col126[93];
   data_col126[95] <= data_col126[94];
   data_col126[96] <= data_col126[95];
   data_col126[97] <= data_col126[96];
   data_col126[98] <= data_col126[97];
   data_col126[99] <= data_col126[98];
   data_col126[100] <= data_col126[99];
   data_col126[101] <= data_col126[100];
   data_col126[102] <= data_col126[101];
   data_col126[103] <= data_col126[102];
   data_col126[104] <= data_col126[103];
   data_col126[105] <= data_col126[104];
   data_col126[106] <= data_col126[105];
   data_col126[107] <= data_col126[106];
   data_col126[108] <= data_col126[107];
   data_col126[109] <= data_col126[108];
   data_col126[110] <= data_col126[109];
   data_col126[111] <= data_col126[110];
   data_col126[112] <= data_col126[111];
   data_col126[113] <= data_col126[112];
   data_col126[114] <= data_col126[113];
   data_col126[115] <= data_col126[114];
   data_col126[116] <= data_col126[115];
   data_col126[117] <= data_col126[116];
   data_col126[118] <= data_col126[117];
   data_col126[119] <= data_col126[118];
   data_col126[120] <= data_col126[119];
   data_col126[121] <= data_col126[120];
   data_col126[122] <= data_col126[121];
   data_col126[123] <= data_col126[122];
   data_col126[124] <= data_col126[123];
   data_col126[125] <= data_col126[124];
   data_col126[126] <= data_col126[125];

   data_col127[1] <= data[38];
   data_col127[2] <= data_col127[1];
   data_col127[3] <= data_col127[2];
   data_col127[4] <= data_col127[3];
   data_col127[5] <= data_col127[4];
   data_col127[6] <= data_col127[5];
   data_col127[7] <= data_col127[6];
   data_col127[8] <= data_col127[7];
   data_col127[9] <= data_col127[8];
   data_col127[10] <= data_col127[9];
   data_col127[11] <= data_col127[10];
   data_col127[12] <= data_col127[11];
   data_col127[13] <= data_col127[12];
   data_col127[14] <= data_col127[13];
   data_col127[15] <= data_col127[14];
   data_col127[16] <= data_col127[15];
   data_col127[17] <= data_col127[16];
   data_col127[18] <= data_col127[17];
   data_col127[19] <= data_col127[18];
   data_col127[20] <= data_col127[19];
   data_col127[21] <= data_col127[20];
   data_col127[22] <= data_col127[21];
   data_col127[23] <= data_col127[22];
   data_col127[24] <= data_col127[23];
   data_col127[25] <= data_col127[24];
   data_col127[26] <= data_col127[25];
   data_col127[27] <= data_col127[26];
   data_col127[28] <= data_col127[27];
   data_col127[29] <= data_col127[28];
   data_col127[30] <= data_col127[29];
   data_col127[31] <= data_col127[30];
   data_col127[32] <= data_col127[31];
   data_col127[33] <= data_col127[32];
   data_col127[34] <= data_col127[33];
   data_col127[35] <= data_col127[34];
   data_col127[36] <= data_col127[35];
   data_col127[37] <= data_col127[36];
   data_col127[38] <= data_col127[37];
   data_col127[39] <= data_col127[38];
   data_col127[40] <= data_col127[39];
   data_col127[41] <= data_col127[40];
   data_col127[42] <= data_col127[41];
   data_col127[43] <= data_col127[42];
   data_col127[44] <= data_col127[43];
   data_col127[45] <= data_col127[44];
   data_col127[46] <= data_col127[45];
   data_col127[47] <= data_col127[46];
   data_col127[48] <= data_col127[47];
   data_col127[49] <= data_col127[48];
   data_col127[50] <= data_col127[49];
   data_col127[51] <= data_col127[50];
   data_col127[52] <= data_col127[51];
   data_col127[53] <= data_col127[52];
   data_col127[54] <= data_col127[53];
   data_col127[55] <= data_col127[54];
   data_col127[56] <= data_col127[55];
   data_col127[57] <= data_col127[56];
   data_col127[58] <= data_col127[57];
   data_col127[59] <= data_col127[58];
   data_col127[60] <= data_col127[59];
   data_col127[61] <= data_col127[60];
   data_col127[62] <= data_col127[61];
   data_col127[63] <= data_col127[62];
   data_col127[64] <= data_col127[63];
   data_col127[65] <= data_col127[64];
   data_col127[66] <= data_col127[65];
   data_col127[67] <= data_col127[66];
   data_col127[68] <= data_col127[67];
   data_col127[69] <= data_col127[68];
   data_col127[70] <= data_col127[69];
   data_col127[71] <= data_col127[70];
   data_col127[72] <= data_col127[71];
   data_col127[73] <= data_col127[72];
   data_col127[74] <= data_col127[73];
   data_col127[75] <= data_col127[74];
   data_col127[76] <= data_col127[75];
   data_col127[77] <= data_col127[76];
   data_col127[78] <= data_col127[77];
   data_col127[79] <= data_col127[78];
   data_col127[80] <= data_col127[79];
   data_col127[81] <= data_col127[80];
   data_col127[82] <= data_col127[81];
   data_col127[83] <= data_col127[82];
   data_col127[84] <= data_col127[83];
   data_col127[85] <= data_col127[84];
   data_col127[86] <= data_col127[85];
   data_col127[87] <= data_col127[86];
   data_col127[88] <= data_col127[87];
   data_col127[89] <= data_col127[88];
   data_col127[90] <= data_col127[89];
   data_col127[91] <= data_col127[90];
   data_col127[92] <= data_col127[91];
   data_col127[93] <= data_col127[92];
   data_col127[94] <= data_col127[93];
   data_col127[95] <= data_col127[94];
   data_col127[96] <= data_col127[95];
   data_col127[97] <= data_col127[96];
   data_col127[98] <= data_col127[97];
   data_col127[99] <= data_col127[98];
   data_col127[100] <= data_col127[99];
   data_col127[101] <= data_col127[100];
   data_col127[102] <= data_col127[101];
   data_col127[103] <= data_col127[102];
   data_col127[104] <= data_col127[103];
   data_col127[105] <= data_col127[104];
   data_col127[106] <= data_col127[105];
   data_col127[107] <= data_col127[106];
   data_col127[108] <= data_col127[107];
   data_col127[109] <= data_col127[108];
   data_col127[110] <= data_col127[109];
   data_col127[111] <= data_col127[110];
   data_col127[112] <= data_col127[111];
   data_col127[113] <= data_col127[112];
   data_col127[114] <= data_col127[113];
   data_col127[115] <= data_col127[114];
   data_col127[116] <= data_col127[115];
   data_col127[117] <= data_col127[116];
   data_col127[118] <= data_col127[117];
   data_col127[119] <= data_col127[118];
   data_col127[120] <= data_col127[119];
   data_col127[121] <= data_col127[120];
   data_col127[122] <= data_col127[121];
   data_col127[123] <= data_col127[122];
   data_col127[124] <= data_col127[123];
   data_col127[125] <= data_col127[124];
   data_col127[126] <= data_col127[125];
   data_col127[127] <= data_col127[126];

   data_col128[1] <= data[37];
   data_col128[2] <= data_col128[1];
   data_col128[3] <= data_col128[2];
   data_col128[4] <= data_col128[3];
   data_col128[5] <= data_col128[4];
   data_col128[6] <= data_col128[5];
   data_col128[7] <= data_col128[6];
   data_col128[8] <= data_col128[7];
   data_col128[9] <= data_col128[8];
   data_col128[10] <= data_col128[9];
   data_col128[11] <= data_col128[10];
   data_col128[12] <= data_col128[11];
   data_col128[13] <= data_col128[12];
   data_col128[14] <= data_col128[13];
   data_col128[15] <= data_col128[14];
   data_col128[16] <= data_col128[15];
   data_col128[17] <= data_col128[16];
   data_col128[18] <= data_col128[17];
   data_col128[19] <= data_col128[18];
   data_col128[20] <= data_col128[19];
   data_col128[21] <= data_col128[20];
   data_col128[22] <= data_col128[21];
   data_col128[23] <= data_col128[22];
   data_col128[24] <= data_col128[23];
   data_col128[25] <= data_col128[24];
   data_col128[26] <= data_col128[25];
   data_col128[27] <= data_col128[26];
   data_col128[28] <= data_col128[27];
   data_col128[29] <= data_col128[28];
   data_col128[30] <= data_col128[29];
   data_col128[31] <= data_col128[30];
   data_col128[32] <= data_col128[31];
   data_col128[33] <= data_col128[32];
   data_col128[34] <= data_col128[33];
   data_col128[35] <= data_col128[34];
   data_col128[36] <= data_col128[35];
   data_col128[37] <= data_col128[36];
   data_col128[38] <= data_col128[37];
   data_col128[39] <= data_col128[38];
   data_col128[40] <= data_col128[39];
   data_col128[41] <= data_col128[40];
   data_col128[42] <= data_col128[41];
   data_col128[43] <= data_col128[42];
   data_col128[44] <= data_col128[43];
   data_col128[45] <= data_col128[44];
   data_col128[46] <= data_col128[45];
   data_col128[47] <= data_col128[46];
   data_col128[48] <= data_col128[47];
   data_col128[49] <= data_col128[48];
   data_col128[50] <= data_col128[49];
   data_col128[51] <= data_col128[50];
   data_col128[52] <= data_col128[51];
   data_col128[53] <= data_col128[52];
   data_col128[54] <= data_col128[53];
   data_col128[55] <= data_col128[54];
   data_col128[56] <= data_col128[55];
   data_col128[57] <= data_col128[56];
   data_col128[58] <= data_col128[57];
   data_col128[59] <= data_col128[58];
   data_col128[60] <= data_col128[59];
   data_col128[61] <= data_col128[60];
   data_col128[62] <= data_col128[61];
   data_col128[63] <= data_col128[62];
   data_col128[64] <= data_col128[63];
   data_col128[65] <= data_col128[64];
   data_col128[66] <= data_col128[65];
   data_col128[67] <= data_col128[66];
   data_col128[68] <= data_col128[67];
   data_col128[69] <= data_col128[68];
   data_col128[70] <= data_col128[69];
   data_col128[71] <= data_col128[70];
   data_col128[72] <= data_col128[71];
   data_col128[73] <= data_col128[72];
   data_col128[74] <= data_col128[73];
   data_col128[75] <= data_col128[74];
   data_col128[76] <= data_col128[75];
   data_col128[77] <= data_col128[76];
   data_col128[78] <= data_col128[77];
   data_col128[79] <= data_col128[78];
   data_col128[80] <= data_col128[79];
   data_col128[81] <= data_col128[80];
   data_col128[82] <= data_col128[81];
   data_col128[83] <= data_col128[82];
   data_col128[84] <= data_col128[83];
   data_col128[85] <= data_col128[84];
   data_col128[86] <= data_col128[85];
   data_col128[87] <= data_col128[86];
   data_col128[88] <= data_col128[87];
   data_col128[89] <= data_col128[88];
   data_col128[90] <= data_col128[89];
   data_col128[91] <= data_col128[90];
   data_col128[92] <= data_col128[91];
   data_col128[93] <= data_col128[92];
   data_col128[94] <= data_col128[93];
   data_col128[95] <= data_col128[94];
   data_col128[96] <= data_col128[95];
   data_col128[97] <= data_col128[96];
   data_col128[98] <= data_col128[97];
   data_col128[99] <= data_col128[98];
   data_col128[100] <= data_col128[99];
   data_col128[101] <= data_col128[100];
   data_col128[102] <= data_col128[101];
   data_col128[103] <= data_col128[102];
   data_col128[104] <= data_col128[103];
   data_col128[105] <= data_col128[104];
   data_col128[106] <= data_col128[105];
   data_col128[107] <= data_col128[106];
   data_col128[108] <= data_col128[107];
   data_col128[109] <= data_col128[108];
   data_col128[110] <= data_col128[109];
   data_col128[111] <= data_col128[110];
   data_col128[112] <= data_col128[111];
   data_col128[113] <= data_col128[112];
   data_col128[114] <= data_col128[113];
   data_col128[115] <= data_col128[114];
   data_col128[116] <= data_col128[115];
   data_col128[117] <= data_col128[116];
   data_col128[118] <= data_col128[117];
   data_col128[119] <= data_col128[118];
   data_col128[120] <= data_col128[119];
   data_col128[121] <= data_col128[120];
   data_col128[122] <= data_col128[121];
   data_col128[123] <= data_col128[122];
   data_col128[124] <= data_col128[123];
   data_col128[125] <= data_col128[124];
   data_col128[126] <= data_col128[125];
   data_col128[127] <= data_col128[126];
   data_col128[128] <= data_col128[127];

   data_col129[1] <= data[36];
   data_col129[2] <= data_col129[1];
   data_col129[3] <= data_col129[2];
   data_col129[4] <= data_col129[3];
   data_col129[5] <= data_col129[4];
   data_col129[6] <= data_col129[5];
   data_col129[7] <= data_col129[6];
   data_col129[8] <= data_col129[7];
   data_col129[9] <= data_col129[8];
   data_col129[10] <= data_col129[9];
   data_col129[11] <= data_col129[10];
   data_col129[12] <= data_col129[11];
   data_col129[13] <= data_col129[12];
   data_col129[14] <= data_col129[13];
   data_col129[15] <= data_col129[14];
   data_col129[16] <= data_col129[15];
   data_col129[17] <= data_col129[16];
   data_col129[18] <= data_col129[17];
   data_col129[19] <= data_col129[18];
   data_col129[20] <= data_col129[19];
   data_col129[21] <= data_col129[20];
   data_col129[22] <= data_col129[21];
   data_col129[23] <= data_col129[22];
   data_col129[24] <= data_col129[23];
   data_col129[25] <= data_col129[24];
   data_col129[26] <= data_col129[25];
   data_col129[27] <= data_col129[26];
   data_col129[28] <= data_col129[27];
   data_col129[29] <= data_col129[28];
   data_col129[30] <= data_col129[29];
   data_col129[31] <= data_col129[30];
   data_col129[32] <= data_col129[31];
   data_col129[33] <= data_col129[32];
   data_col129[34] <= data_col129[33];
   data_col129[35] <= data_col129[34];
   data_col129[36] <= data_col129[35];
   data_col129[37] <= data_col129[36];
   data_col129[38] <= data_col129[37];
   data_col129[39] <= data_col129[38];
   data_col129[40] <= data_col129[39];
   data_col129[41] <= data_col129[40];
   data_col129[42] <= data_col129[41];
   data_col129[43] <= data_col129[42];
   data_col129[44] <= data_col129[43];
   data_col129[45] <= data_col129[44];
   data_col129[46] <= data_col129[45];
   data_col129[47] <= data_col129[46];
   data_col129[48] <= data_col129[47];
   data_col129[49] <= data_col129[48];
   data_col129[50] <= data_col129[49];
   data_col129[51] <= data_col129[50];
   data_col129[52] <= data_col129[51];
   data_col129[53] <= data_col129[52];
   data_col129[54] <= data_col129[53];
   data_col129[55] <= data_col129[54];
   data_col129[56] <= data_col129[55];
   data_col129[57] <= data_col129[56];
   data_col129[58] <= data_col129[57];
   data_col129[59] <= data_col129[58];
   data_col129[60] <= data_col129[59];
   data_col129[61] <= data_col129[60];
   data_col129[62] <= data_col129[61];
   data_col129[63] <= data_col129[62];
   data_col129[64] <= data_col129[63];
   data_col129[65] <= data_col129[64];
   data_col129[66] <= data_col129[65];
   data_col129[67] <= data_col129[66];
   data_col129[68] <= data_col129[67];
   data_col129[69] <= data_col129[68];
   data_col129[70] <= data_col129[69];
   data_col129[71] <= data_col129[70];
   data_col129[72] <= data_col129[71];
   data_col129[73] <= data_col129[72];
   data_col129[74] <= data_col129[73];
   data_col129[75] <= data_col129[74];
   data_col129[76] <= data_col129[75];
   data_col129[77] <= data_col129[76];
   data_col129[78] <= data_col129[77];
   data_col129[79] <= data_col129[78];
   data_col129[80] <= data_col129[79];
   data_col129[81] <= data_col129[80];
   data_col129[82] <= data_col129[81];
   data_col129[83] <= data_col129[82];
   data_col129[84] <= data_col129[83];
   data_col129[85] <= data_col129[84];
   data_col129[86] <= data_col129[85];
   data_col129[87] <= data_col129[86];
   data_col129[88] <= data_col129[87];
   data_col129[89] <= data_col129[88];
   data_col129[90] <= data_col129[89];
   data_col129[91] <= data_col129[90];
   data_col129[92] <= data_col129[91];
   data_col129[93] <= data_col129[92];
   data_col129[94] <= data_col129[93];
   data_col129[95] <= data_col129[94];
   data_col129[96] <= data_col129[95];
   data_col129[97] <= data_col129[96];
   data_col129[98] <= data_col129[97];
   data_col129[99] <= data_col129[98];
   data_col129[100] <= data_col129[99];
   data_col129[101] <= data_col129[100];
   data_col129[102] <= data_col129[101];
   data_col129[103] <= data_col129[102];
   data_col129[104] <= data_col129[103];
   data_col129[105] <= data_col129[104];
   data_col129[106] <= data_col129[105];
   data_col129[107] <= data_col129[106];
   data_col129[108] <= data_col129[107];
   data_col129[109] <= data_col129[108];
   data_col129[110] <= data_col129[109];
   data_col129[111] <= data_col129[110];
   data_col129[112] <= data_col129[111];
   data_col129[113] <= data_col129[112];
   data_col129[114] <= data_col129[113];
   data_col129[115] <= data_col129[114];
   data_col129[116] <= data_col129[115];
   data_col129[117] <= data_col129[116];
   data_col129[118] <= data_col129[117];
   data_col129[119] <= data_col129[118];
   data_col129[120] <= data_col129[119];
   data_col129[121] <= data_col129[120];
   data_col129[122] <= data_col129[121];
   data_col129[123] <= data_col129[122];
   data_col129[124] <= data_col129[123];
   data_col129[125] <= data_col129[124];
   data_col129[126] <= data_col129[125];
   data_col129[127] <= data_col129[126];
   data_col129[128] <= data_col129[127];
   data_col129[129] <= data_col129[128];

   data_col130[1] <= data[35];
   data_col130[2] <= data_col130[1];
   data_col130[3] <= data_col130[2];
   data_col130[4] <= data_col130[3];
   data_col130[5] <= data_col130[4];
   data_col130[6] <= data_col130[5];
   data_col130[7] <= data_col130[6];
   data_col130[8] <= data_col130[7];
   data_col130[9] <= data_col130[8];
   data_col130[10] <= data_col130[9];
   data_col130[11] <= data_col130[10];
   data_col130[12] <= data_col130[11];
   data_col130[13] <= data_col130[12];
   data_col130[14] <= data_col130[13];
   data_col130[15] <= data_col130[14];
   data_col130[16] <= data_col130[15];
   data_col130[17] <= data_col130[16];
   data_col130[18] <= data_col130[17];
   data_col130[19] <= data_col130[18];
   data_col130[20] <= data_col130[19];
   data_col130[21] <= data_col130[20];
   data_col130[22] <= data_col130[21];
   data_col130[23] <= data_col130[22];
   data_col130[24] <= data_col130[23];
   data_col130[25] <= data_col130[24];
   data_col130[26] <= data_col130[25];
   data_col130[27] <= data_col130[26];
   data_col130[28] <= data_col130[27];
   data_col130[29] <= data_col130[28];
   data_col130[30] <= data_col130[29];
   data_col130[31] <= data_col130[30];
   data_col130[32] <= data_col130[31];
   data_col130[33] <= data_col130[32];
   data_col130[34] <= data_col130[33];
   data_col130[35] <= data_col130[34];
   data_col130[36] <= data_col130[35];
   data_col130[37] <= data_col130[36];
   data_col130[38] <= data_col130[37];
   data_col130[39] <= data_col130[38];
   data_col130[40] <= data_col130[39];
   data_col130[41] <= data_col130[40];
   data_col130[42] <= data_col130[41];
   data_col130[43] <= data_col130[42];
   data_col130[44] <= data_col130[43];
   data_col130[45] <= data_col130[44];
   data_col130[46] <= data_col130[45];
   data_col130[47] <= data_col130[46];
   data_col130[48] <= data_col130[47];
   data_col130[49] <= data_col130[48];
   data_col130[50] <= data_col130[49];
   data_col130[51] <= data_col130[50];
   data_col130[52] <= data_col130[51];
   data_col130[53] <= data_col130[52];
   data_col130[54] <= data_col130[53];
   data_col130[55] <= data_col130[54];
   data_col130[56] <= data_col130[55];
   data_col130[57] <= data_col130[56];
   data_col130[58] <= data_col130[57];
   data_col130[59] <= data_col130[58];
   data_col130[60] <= data_col130[59];
   data_col130[61] <= data_col130[60];
   data_col130[62] <= data_col130[61];
   data_col130[63] <= data_col130[62];
   data_col130[64] <= data_col130[63];
   data_col130[65] <= data_col130[64];
   data_col130[66] <= data_col130[65];
   data_col130[67] <= data_col130[66];
   data_col130[68] <= data_col130[67];
   data_col130[69] <= data_col130[68];
   data_col130[70] <= data_col130[69];
   data_col130[71] <= data_col130[70];
   data_col130[72] <= data_col130[71];
   data_col130[73] <= data_col130[72];
   data_col130[74] <= data_col130[73];
   data_col130[75] <= data_col130[74];
   data_col130[76] <= data_col130[75];
   data_col130[77] <= data_col130[76];
   data_col130[78] <= data_col130[77];
   data_col130[79] <= data_col130[78];
   data_col130[80] <= data_col130[79];
   data_col130[81] <= data_col130[80];
   data_col130[82] <= data_col130[81];
   data_col130[83] <= data_col130[82];
   data_col130[84] <= data_col130[83];
   data_col130[85] <= data_col130[84];
   data_col130[86] <= data_col130[85];
   data_col130[87] <= data_col130[86];
   data_col130[88] <= data_col130[87];
   data_col130[89] <= data_col130[88];
   data_col130[90] <= data_col130[89];
   data_col130[91] <= data_col130[90];
   data_col130[92] <= data_col130[91];
   data_col130[93] <= data_col130[92];
   data_col130[94] <= data_col130[93];
   data_col130[95] <= data_col130[94];
   data_col130[96] <= data_col130[95];
   data_col130[97] <= data_col130[96];
   data_col130[98] <= data_col130[97];
   data_col130[99] <= data_col130[98];
   data_col130[100] <= data_col130[99];
   data_col130[101] <= data_col130[100];
   data_col130[102] <= data_col130[101];
   data_col130[103] <= data_col130[102];
   data_col130[104] <= data_col130[103];
   data_col130[105] <= data_col130[104];
   data_col130[106] <= data_col130[105];
   data_col130[107] <= data_col130[106];
   data_col130[108] <= data_col130[107];
   data_col130[109] <= data_col130[108];
   data_col130[110] <= data_col130[109];
   data_col130[111] <= data_col130[110];
   data_col130[112] <= data_col130[111];
   data_col130[113] <= data_col130[112];
   data_col130[114] <= data_col130[113];
   data_col130[115] <= data_col130[114];
   data_col130[116] <= data_col130[115];
   data_col130[117] <= data_col130[116];
   data_col130[118] <= data_col130[117];
   data_col130[119] <= data_col130[118];
   data_col130[120] <= data_col130[119];
   data_col130[121] <= data_col130[120];
   data_col130[122] <= data_col130[121];
   data_col130[123] <= data_col130[122];
   data_col130[124] <= data_col130[123];
   data_col130[125] <= data_col130[124];
   data_col130[126] <= data_col130[125];
   data_col130[127] <= data_col130[126];
   data_col130[128] <= data_col130[127];
   data_col130[129] <= data_col130[128];
   data_col130[130] <= data_col130[129];

   data_col131[1] <= data[34];
   data_col131[2] <= data_col131[1];
   data_col131[3] <= data_col131[2];
   data_col131[4] <= data_col131[3];
   data_col131[5] <= data_col131[4];
   data_col131[6] <= data_col131[5];
   data_col131[7] <= data_col131[6];
   data_col131[8] <= data_col131[7];
   data_col131[9] <= data_col131[8];
   data_col131[10] <= data_col131[9];
   data_col131[11] <= data_col131[10];
   data_col131[12] <= data_col131[11];
   data_col131[13] <= data_col131[12];
   data_col131[14] <= data_col131[13];
   data_col131[15] <= data_col131[14];
   data_col131[16] <= data_col131[15];
   data_col131[17] <= data_col131[16];
   data_col131[18] <= data_col131[17];
   data_col131[19] <= data_col131[18];
   data_col131[20] <= data_col131[19];
   data_col131[21] <= data_col131[20];
   data_col131[22] <= data_col131[21];
   data_col131[23] <= data_col131[22];
   data_col131[24] <= data_col131[23];
   data_col131[25] <= data_col131[24];
   data_col131[26] <= data_col131[25];
   data_col131[27] <= data_col131[26];
   data_col131[28] <= data_col131[27];
   data_col131[29] <= data_col131[28];
   data_col131[30] <= data_col131[29];
   data_col131[31] <= data_col131[30];
   data_col131[32] <= data_col131[31];
   data_col131[33] <= data_col131[32];
   data_col131[34] <= data_col131[33];
   data_col131[35] <= data_col131[34];
   data_col131[36] <= data_col131[35];
   data_col131[37] <= data_col131[36];
   data_col131[38] <= data_col131[37];
   data_col131[39] <= data_col131[38];
   data_col131[40] <= data_col131[39];
   data_col131[41] <= data_col131[40];
   data_col131[42] <= data_col131[41];
   data_col131[43] <= data_col131[42];
   data_col131[44] <= data_col131[43];
   data_col131[45] <= data_col131[44];
   data_col131[46] <= data_col131[45];
   data_col131[47] <= data_col131[46];
   data_col131[48] <= data_col131[47];
   data_col131[49] <= data_col131[48];
   data_col131[50] <= data_col131[49];
   data_col131[51] <= data_col131[50];
   data_col131[52] <= data_col131[51];
   data_col131[53] <= data_col131[52];
   data_col131[54] <= data_col131[53];
   data_col131[55] <= data_col131[54];
   data_col131[56] <= data_col131[55];
   data_col131[57] <= data_col131[56];
   data_col131[58] <= data_col131[57];
   data_col131[59] <= data_col131[58];
   data_col131[60] <= data_col131[59];
   data_col131[61] <= data_col131[60];
   data_col131[62] <= data_col131[61];
   data_col131[63] <= data_col131[62];
   data_col131[64] <= data_col131[63];
   data_col131[65] <= data_col131[64];
   data_col131[66] <= data_col131[65];
   data_col131[67] <= data_col131[66];
   data_col131[68] <= data_col131[67];
   data_col131[69] <= data_col131[68];
   data_col131[70] <= data_col131[69];
   data_col131[71] <= data_col131[70];
   data_col131[72] <= data_col131[71];
   data_col131[73] <= data_col131[72];
   data_col131[74] <= data_col131[73];
   data_col131[75] <= data_col131[74];
   data_col131[76] <= data_col131[75];
   data_col131[77] <= data_col131[76];
   data_col131[78] <= data_col131[77];
   data_col131[79] <= data_col131[78];
   data_col131[80] <= data_col131[79];
   data_col131[81] <= data_col131[80];
   data_col131[82] <= data_col131[81];
   data_col131[83] <= data_col131[82];
   data_col131[84] <= data_col131[83];
   data_col131[85] <= data_col131[84];
   data_col131[86] <= data_col131[85];
   data_col131[87] <= data_col131[86];
   data_col131[88] <= data_col131[87];
   data_col131[89] <= data_col131[88];
   data_col131[90] <= data_col131[89];
   data_col131[91] <= data_col131[90];
   data_col131[92] <= data_col131[91];
   data_col131[93] <= data_col131[92];
   data_col131[94] <= data_col131[93];
   data_col131[95] <= data_col131[94];
   data_col131[96] <= data_col131[95];
   data_col131[97] <= data_col131[96];
   data_col131[98] <= data_col131[97];
   data_col131[99] <= data_col131[98];
   data_col131[100] <= data_col131[99];
   data_col131[101] <= data_col131[100];
   data_col131[102] <= data_col131[101];
   data_col131[103] <= data_col131[102];
   data_col131[104] <= data_col131[103];
   data_col131[105] <= data_col131[104];
   data_col131[106] <= data_col131[105];
   data_col131[107] <= data_col131[106];
   data_col131[108] <= data_col131[107];
   data_col131[109] <= data_col131[108];
   data_col131[110] <= data_col131[109];
   data_col131[111] <= data_col131[110];
   data_col131[112] <= data_col131[111];
   data_col131[113] <= data_col131[112];
   data_col131[114] <= data_col131[113];
   data_col131[115] <= data_col131[114];
   data_col131[116] <= data_col131[115];
   data_col131[117] <= data_col131[116];
   data_col131[118] <= data_col131[117];
   data_col131[119] <= data_col131[118];
   data_col131[120] <= data_col131[119];
   data_col131[121] <= data_col131[120];
   data_col131[122] <= data_col131[121];
   data_col131[123] <= data_col131[122];
   data_col131[124] <= data_col131[123];
   data_col131[125] <= data_col131[124];
   data_col131[126] <= data_col131[125];
   data_col131[127] <= data_col131[126];
   data_col131[128] <= data_col131[127];
   data_col131[129] <= data_col131[128];
   data_col131[130] <= data_col131[129];
   data_col131[131] <= data_col131[130];

   data_col132[1] <= data[33];
   data_col132[2] <= data_col132[1];
   data_col132[3] <= data_col132[2];
   data_col132[4] <= data_col132[3];
   data_col132[5] <= data_col132[4];
   data_col132[6] <= data_col132[5];
   data_col132[7] <= data_col132[6];
   data_col132[8] <= data_col132[7];
   data_col132[9] <= data_col132[8];
   data_col132[10] <= data_col132[9];
   data_col132[11] <= data_col132[10];
   data_col132[12] <= data_col132[11];
   data_col132[13] <= data_col132[12];
   data_col132[14] <= data_col132[13];
   data_col132[15] <= data_col132[14];
   data_col132[16] <= data_col132[15];
   data_col132[17] <= data_col132[16];
   data_col132[18] <= data_col132[17];
   data_col132[19] <= data_col132[18];
   data_col132[20] <= data_col132[19];
   data_col132[21] <= data_col132[20];
   data_col132[22] <= data_col132[21];
   data_col132[23] <= data_col132[22];
   data_col132[24] <= data_col132[23];
   data_col132[25] <= data_col132[24];
   data_col132[26] <= data_col132[25];
   data_col132[27] <= data_col132[26];
   data_col132[28] <= data_col132[27];
   data_col132[29] <= data_col132[28];
   data_col132[30] <= data_col132[29];
   data_col132[31] <= data_col132[30];
   data_col132[32] <= data_col132[31];
   data_col132[33] <= data_col132[32];
   data_col132[34] <= data_col132[33];
   data_col132[35] <= data_col132[34];
   data_col132[36] <= data_col132[35];
   data_col132[37] <= data_col132[36];
   data_col132[38] <= data_col132[37];
   data_col132[39] <= data_col132[38];
   data_col132[40] <= data_col132[39];
   data_col132[41] <= data_col132[40];
   data_col132[42] <= data_col132[41];
   data_col132[43] <= data_col132[42];
   data_col132[44] <= data_col132[43];
   data_col132[45] <= data_col132[44];
   data_col132[46] <= data_col132[45];
   data_col132[47] <= data_col132[46];
   data_col132[48] <= data_col132[47];
   data_col132[49] <= data_col132[48];
   data_col132[50] <= data_col132[49];
   data_col132[51] <= data_col132[50];
   data_col132[52] <= data_col132[51];
   data_col132[53] <= data_col132[52];
   data_col132[54] <= data_col132[53];
   data_col132[55] <= data_col132[54];
   data_col132[56] <= data_col132[55];
   data_col132[57] <= data_col132[56];
   data_col132[58] <= data_col132[57];
   data_col132[59] <= data_col132[58];
   data_col132[60] <= data_col132[59];
   data_col132[61] <= data_col132[60];
   data_col132[62] <= data_col132[61];
   data_col132[63] <= data_col132[62];
   data_col132[64] <= data_col132[63];
   data_col132[65] <= data_col132[64];
   data_col132[66] <= data_col132[65];
   data_col132[67] <= data_col132[66];
   data_col132[68] <= data_col132[67];
   data_col132[69] <= data_col132[68];
   data_col132[70] <= data_col132[69];
   data_col132[71] <= data_col132[70];
   data_col132[72] <= data_col132[71];
   data_col132[73] <= data_col132[72];
   data_col132[74] <= data_col132[73];
   data_col132[75] <= data_col132[74];
   data_col132[76] <= data_col132[75];
   data_col132[77] <= data_col132[76];
   data_col132[78] <= data_col132[77];
   data_col132[79] <= data_col132[78];
   data_col132[80] <= data_col132[79];
   data_col132[81] <= data_col132[80];
   data_col132[82] <= data_col132[81];
   data_col132[83] <= data_col132[82];
   data_col132[84] <= data_col132[83];
   data_col132[85] <= data_col132[84];
   data_col132[86] <= data_col132[85];
   data_col132[87] <= data_col132[86];
   data_col132[88] <= data_col132[87];
   data_col132[89] <= data_col132[88];
   data_col132[90] <= data_col132[89];
   data_col132[91] <= data_col132[90];
   data_col132[92] <= data_col132[91];
   data_col132[93] <= data_col132[92];
   data_col132[94] <= data_col132[93];
   data_col132[95] <= data_col132[94];
   data_col132[96] <= data_col132[95];
   data_col132[97] <= data_col132[96];
   data_col132[98] <= data_col132[97];
   data_col132[99] <= data_col132[98];
   data_col132[100] <= data_col132[99];
   data_col132[101] <= data_col132[100];
   data_col132[102] <= data_col132[101];
   data_col132[103] <= data_col132[102];
   data_col132[104] <= data_col132[103];
   data_col132[105] <= data_col132[104];
   data_col132[106] <= data_col132[105];
   data_col132[107] <= data_col132[106];
   data_col132[108] <= data_col132[107];
   data_col132[109] <= data_col132[108];
   data_col132[110] <= data_col132[109];
   data_col132[111] <= data_col132[110];
   data_col132[112] <= data_col132[111];
   data_col132[113] <= data_col132[112];
   data_col132[114] <= data_col132[113];
   data_col132[115] <= data_col132[114];
   data_col132[116] <= data_col132[115];
   data_col132[117] <= data_col132[116];
   data_col132[118] <= data_col132[117];
   data_col132[119] <= data_col132[118];
   data_col132[120] <= data_col132[119];
   data_col132[121] <= data_col132[120];
   data_col132[122] <= data_col132[121];
   data_col132[123] <= data_col132[122];
   data_col132[124] <= data_col132[123];
   data_col132[125] <= data_col132[124];
   data_col132[126] <= data_col132[125];
   data_col132[127] <= data_col132[126];
   data_col132[128] <= data_col132[127];
   data_col132[129] <= data_col132[128];
   data_col132[130] <= data_col132[129];
   data_col132[131] <= data_col132[130];
   data_col132[132] <= data_col132[131];

   data_col133[1] <= data[32];
   data_col133[2] <= data_col133[1];
   data_col133[3] <= data_col133[2];
   data_col133[4] <= data_col133[3];
   data_col133[5] <= data_col133[4];
   data_col133[6] <= data_col133[5];
   data_col133[7] <= data_col133[6];
   data_col133[8] <= data_col133[7];
   data_col133[9] <= data_col133[8];
   data_col133[10] <= data_col133[9];
   data_col133[11] <= data_col133[10];
   data_col133[12] <= data_col133[11];
   data_col133[13] <= data_col133[12];
   data_col133[14] <= data_col133[13];
   data_col133[15] <= data_col133[14];
   data_col133[16] <= data_col133[15];
   data_col133[17] <= data_col133[16];
   data_col133[18] <= data_col133[17];
   data_col133[19] <= data_col133[18];
   data_col133[20] <= data_col133[19];
   data_col133[21] <= data_col133[20];
   data_col133[22] <= data_col133[21];
   data_col133[23] <= data_col133[22];
   data_col133[24] <= data_col133[23];
   data_col133[25] <= data_col133[24];
   data_col133[26] <= data_col133[25];
   data_col133[27] <= data_col133[26];
   data_col133[28] <= data_col133[27];
   data_col133[29] <= data_col133[28];
   data_col133[30] <= data_col133[29];
   data_col133[31] <= data_col133[30];
   data_col133[32] <= data_col133[31];
   data_col133[33] <= data_col133[32];
   data_col133[34] <= data_col133[33];
   data_col133[35] <= data_col133[34];
   data_col133[36] <= data_col133[35];
   data_col133[37] <= data_col133[36];
   data_col133[38] <= data_col133[37];
   data_col133[39] <= data_col133[38];
   data_col133[40] <= data_col133[39];
   data_col133[41] <= data_col133[40];
   data_col133[42] <= data_col133[41];
   data_col133[43] <= data_col133[42];
   data_col133[44] <= data_col133[43];
   data_col133[45] <= data_col133[44];
   data_col133[46] <= data_col133[45];
   data_col133[47] <= data_col133[46];
   data_col133[48] <= data_col133[47];
   data_col133[49] <= data_col133[48];
   data_col133[50] <= data_col133[49];
   data_col133[51] <= data_col133[50];
   data_col133[52] <= data_col133[51];
   data_col133[53] <= data_col133[52];
   data_col133[54] <= data_col133[53];
   data_col133[55] <= data_col133[54];
   data_col133[56] <= data_col133[55];
   data_col133[57] <= data_col133[56];
   data_col133[58] <= data_col133[57];
   data_col133[59] <= data_col133[58];
   data_col133[60] <= data_col133[59];
   data_col133[61] <= data_col133[60];
   data_col133[62] <= data_col133[61];
   data_col133[63] <= data_col133[62];
   data_col133[64] <= data_col133[63];
   data_col133[65] <= data_col133[64];
   data_col133[66] <= data_col133[65];
   data_col133[67] <= data_col133[66];
   data_col133[68] <= data_col133[67];
   data_col133[69] <= data_col133[68];
   data_col133[70] <= data_col133[69];
   data_col133[71] <= data_col133[70];
   data_col133[72] <= data_col133[71];
   data_col133[73] <= data_col133[72];
   data_col133[74] <= data_col133[73];
   data_col133[75] <= data_col133[74];
   data_col133[76] <= data_col133[75];
   data_col133[77] <= data_col133[76];
   data_col133[78] <= data_col133[77];
   data_col133[79] <= data_col133[78];
   data_col133[80] <= data_col133[79];
   data_col133[81] <= data_col133[80];
   data_col133[82] <= data_col133[81];
   data_col133[83] <= data_col133[82];
   data_col133[84] <= data_col133[83];
   data_col133[85] <= data_col133[84];
   data_col133[86] <= data_col133[85];
   data_col133[87] <= data_col133[86];
   data_col133[88] <= data_col133[87];
   data_col133[89] <= data_col133[88];
   data_col133[90] <= data_col133[89];
   data_col133[91] <= data_col133[90];
   data_col133[92] <= data_col133[91];
   data_col133[93] <= data_col133[92];
   data_col133[94] <= data_col133[93];
   data_col133[95] <= data_col133[94];
   data_col133[96] <= data_col133[95];
   data_col133[97] <= data_col133[96];
   data_col133[98] <= data_col133[97];
   data_col133[99] <= data_col133[98];
   data_col133[100] <= data_col133[99];
   data_col133[101] <= data_col133[100];
   data_col133[102] <= data_col133[101];
   data_col133[103] <= data_col133[102];
   data_col133[104] <= data_col133[103];
   data_col133[105] <= data_col133[104];
   data_col133[106] <= data_col133[105];
   data_col133[107] <= data_col133[106];
   data_col133[108] <= data_col133[107];
   data_col133[109] <= data_col133[108];
   data_col133[110] <= data_col133[109];
   data_col133[111] <= data_col133[110];
   data_col133[112] <= data_col133[111];
   data_col133[113] <= data_col133[112];
   data_col133[114] <= data_col133[113];
   data_col133[115] <= data_col133[114];
   data_col133[116] <= data_col133[115];
   data_col133[117] <= data_col133[116];
   data_col133[118] <= data_col133[117];
   data_col133[119] <= data_col133[118];
   data_col133[120] <= data_col133[119];
   data_col133[121] <= data_col133[120];
   data_col133[122] <= data_col133[121];
   data_col133[123] <= data_col133[122];
   data_col133[124] <= data_col133[123];
   data_col133[125] <= data_col133[124];
   data_col133[126] <= data_col133[125];
   data_col133[127] <= data_col133[126];
   data_col133[128] <= data_col133[127];
   data_col133[129] <= data_col133[128];
   data_col133[130] <= data_col133[129];
   data_col133[131] <= data_col133[130];
   data_col133[132] <= data_col133[131];
   data_col133[133] <= data_col133[132];

   data_col134[1] <= data[31];
   data_col134[2] <= data_col134[1];
   data_col134[3] <= data_col134[2];
   data_col134[4] <= data_col134[3];
   data_col134[5] <= data_col134[4];
   data_col134[6] <= data_col134[5];
   data_col134[7] <= data_col134[6];
   data_col134[8] <= data_col134[7];
   data_col134[9] <= data_col134[8];
   data_col134[10] <= data_col134[9];
   data_col134[11] <= data_col134[10];
   data_col134[12] <= data_col134[11];
   data_col134[13] <= data_col134[12];
   data_col134[14] <= data_col134[13];
   data_col134[15] <= data_col134[14];
   data_col134[16] <= data_col134[15];
   data_col134[17] <= data_col134[16];
   data_col134[18] <= data_col134[17];
   data_col134[19] <= data_col134[18];
   data_col134[20] <= data_col134[19];
   data_col134[21] <= data_col134[20];
   data_col134[22] <= data_col134[21];
   data_col134[23] <= data_col134[22];
   data_col134[24] <= data_col134[23];
   data_col134[25] <= data_col134[24];
   data_col134[26] <= data_col134[25];
   data_col134[27] <= data_col134[26];
   data_col134[28] <= data_col134[27];
   data_col134[29] <= data_col134[28];
   data_col134[30] <= data_col134[29];
   data_col134[31] <= data_col134[30];
   data_col134[32] <= data_col134[31];
   data_col134[33] <= data_col134[32];
   data_col134[34] <= data_col134[33];
   data_col134[35] <= data_col134[34];
   data_col134[36] <= data_col134[35];
   data_col134[37] <= data_col134[36];
   data_col134[38] <= data_col134[37];
   data_col134[39] <= data_col134[38];
   data_col134[40] <= data_col134[39];
   data_col134[41] <= data_col134[40];
   data_col134[42] <= data_col134[41];
   data_col134[43] <= data_col134[42];
   data_col134[44] <= data_col134[43];
   data_col134[45] <= data_col134[44];
   data_col134[46] <= data_col134[45];
   data_col134[47] <= data_col134[46];
   data_col134[48] <= data_col134[47];
   data_col134[49] <= data_col134[48];
   data_col134[50] <= data_col134[49];
   data_col134[51] <= data_col134[50];
   data_col134[52] <= data_col134[51];
   data_col134[53] <= data_col134[52];
   data_col134[54] <= data_col134[53];
   data_col134[55] <= data_col134[54];
   data_col134[56] <= data_col134[55];
   data_col134[57] <= data_col134[56];
   data_col134[58] <= data_col134[57];
   data_col134[59] <= data_col134[58];
   data_col134[60] <= data_col134[59];
   data_col134[61] <= data_col134[60];
   data_col134[62] <= data_col134[61];
   data_col134[63] <= data_col134[62];
   data_col134[64] <= data_col134[63];
   data_col134[65] <= data_col134[64];
   data_col134[66] <= data_col134[65];
   data_col134[67] <= data_col134[66];
   data_col134[68] <= data_col134[67];
   data_col134[69] <= data_col134[68];
   data_col134[70] <= data_col134[69];
   data_col134[71] <= data_col134[70];
   data_col134[72] <= data_col134[71];
   data_col134[73] <= data_col134[72];
   data_col134[74] <= data_col134[73];
   data_col134[75] <= data_col134[74];
   data_col134[76] <= data_col134[75];
   data_col134[77] <= data_col134[76];
   data_col134[78] <= data_col134[77];
   data_col134[79] <= data_col134[78];
   data_col134[80] <= data_col134[79];
   data_col134[81] <= data_col134[80];
   data_col134[82] <= data_col134[81];
   data_col134[83] <= data_col134[82];
   data_col134[84] <= data_col134[83];
   data_col134[85] <= data_col134[84];
   data_col134[86] <= data_col134[85];
   data_col134[87] <= data_col134[86];
   data_col134[88] <= data_col134[87];
   data_col134[89] <= data_col134[88];
   data_col134[90] <= data_col134[89];
   data_col134[91] <= data_col134[90];
   data_col134[92] <= data_col134[91];
   data_col134[93] <= data_col134[92];
   data_col134[94] <= data_col134[93];
   data_col134[95] <= data_col134[94];
   data_col134[96] <= data_col134[95];
   data_col134[97] <= data_col134[96];
   data_col134[98] <= data_col134[97];
   data_col134[99] <= data_col134[98];
   data_col134[100] <= data_col134[99];
   data_col134[101] <= data_col134[100];
   data_col134[102] <= data_col134[101];
   data_col134[103] <= data_col134[102];
   data_col134[104] <= data_col134[103];
   data_col134[105] <= data_col134[104];
   data_col134[106] <= data_col134[105];
   data_col134[107] <= data_col134[106];
   data_col134[108] <= data_col134[107];
   data_col134[109] <= data_col134[108];
   data_col134[110] <= data_col134[109];
   data_col134[111] <= data_col134[110];
   data_col134[112] <= data_col134[111];
   data_col134[113] <= data_col134[112];
   data_col134[114] <= data_col134[113];
   data_col134[115] <= data_col134[114];
   data_col134[116] <= data_col134[115];
   data_col134[117] <= data_col134[116];
   data_col134[118] <= data_col134[117];
   data_col134[119] <= data_col134[118];
   data_col134[120] <= data_col134[119];
   data_col134[121] <= data_col134[120];
   data_col134[122] <= data_col134[121];
   data_col134[123] <= data_col134[122];
   data_col134[124] <= data_col134[123];
   data_col134[125] <= data_col134[124];
   data_col134[126] <= data_col134[125];
   data_col134[127] <= data_col134[126];
   data_col134[128] <= data_col134[127];
   data_col134[129] <= data_col134[128];
   data_col134[130] <= data_col134[129];
   data_col134[131] <= data_col134[130];
   data_col134[132] <= data_col134[131];
   data_col134[133] <= data_col134[132];
   data_col134[134] <= data_col134[133];

   data_col135[1] <= data[30];
   data_col135[2] <= data_col135[1];
   data_col135[3] <= data_col135[2];
   data_col135[4] <= data_col135[3];
   data_col135[5] <= data_col135[4];
   data_col135[6] <= data_col135[5];
   data_col135[7] <= data_col135[6];
   data_col135[8] <= data_col135[7];
   data_col135[9] <= data_col135[8];
   data_col135[10] <= data_col135[9];
   data_col135[11] <= data_col135[10];
   data_col135[12] <= data_col135[11];
   data_col135[13] <= data_col135[12];
   data_col135[14] <= data_col135[13];
   data_col135[15] <= data_col135[14];
   data_col135[16] <= data_col135[15];
   data_col135[17] <= data_col135[16];
   data_col135[18] <= data_col135[17];
   data_col135[19] <= data_col135[18];
   data_col135[20] <= data_col135[19];
   data_col135[21] <= data_col135[20];
   data_col135[22] <= data_col135[21];
   data_col135[23] <= data_col135[22];
   data_col135[24] <= data_col135[23];
   data_col135[25] <= data_col135[24];
   data_col135[26] <= data_col135[25];
   data_col135[27] <= data_col135[26];
   data_col135[28] <= data_col135[27];
   data_col135[29] <= data_col135[28];
   data_col135[30] <= data_col135[29];
   data_col135[31] <= data_col135[30];
   data_col135[32] <= data_col135[31];
   data_col135[33] <= data_col135[32];
   data_col135[34] <= data_col135[33];
   data_col135[35] <= data_col135[34];
   data_col135[36] <= data_col135[35];
   data_col135[37] <= data_col135[36];
   data_col135[38] <= data_col135[37];
   data_col135[39] <= data_col135[38];
   data_col135[40] <= data_col135[39];
   data_col135[41] <= data_col135[40];
   data_col135[42] <= data_col135[41];
   data_col135[43] <= data_col135[42];
   data_col135[44] <= data_col135[43];
   data_col135[45] <= data_col135[44];
   data_col135[46] <= data_col135[45];
   data_col135[47] <= data_col135[46];
   data_col135[48] <= data_col135[47];
   data_col135[49] <= data_col135[48];
   data_col135[50] <= data_col135[49];
   data_col135[51] <= data_col135[50];
   data_col135[52] <= data_col135[51];
   data_col135[53] <= data_col135[52];
   data_col135[54] <= data_col135[53];
   data_col135[55] <= data_col135[54];
   data_col135[56] <= data_col135[55];
   data_col135[57] <= data_col135[56];
   data_col135[58] <= data_col135[57];
   data_col135[59] <= data_col135[58];
   data_col135[60] <= data_col135[59];
   data_col135[61] <= data_col135[60];
   data_col135[62] <= data_col135[61];
   data_col135[63] <= data_col135[62];
   data_col135[64] <= data_col135[63];
   data_col135[65] <= data_col135[64];
   data_col135[66] <= data_col135[65];
   data_col135[67] <= data_col135[66];
   data_col135[68] <= data_col135[67];
   data_col135[69] <= data_col135[68];
   data_col135[70] <= data_col135[69];
   data_col135[71] <= data_col135[70];
   data_col135[72] <= data_col135[71];
   data_col135[73] <= data_col135[72];
   data_col135[74] <= data_col135[73];
   data_col135[75] <= data_col135[74];
   data_col135[76] <= data_col135[75];
   data_col135[77] <= data_col135[76];
   data_col135[78] <= data_col135[77];
   data_col135[79] <= data_col135[78];
   data_col135[80] <= data_col135[79];
   data_col135[81] <= data_col135[80];
   data_col135[82] <= data_col135[81];
   data_col135[83] <= data_col135[82];
   data_col135[84] <= data_col135[83];
   data_col135[85] <= data_col135[84];
   data_col135[86] <= data_col135[85];
   data_col135[87] <= data_col135[86];
   data_col135[88] <= data_col135[87];
   data_col135[89] <= data_col135[88];
   data_col135[90] <= data_col135[89];
   data_col135[91] <= data_col135[90];
   data_col135[92] <= data_col135[91];
   data_col135[93] <= data_col135[92];
   data_col135[94] <= data_col135[93];
   data_col135[95] <= data_col135[94];
   data_col135[96] <= data_col135[95];
   data_col135[97] <= data_col135[96];
   data_col135[98] <= data_col135[97];
   data_col135[99] <= data_col135[98];
   data_col135[100] <= data_col135[99];
   data_col135[101] <= data_col135[100];
   data_col135[102] <= data_col135[101];
   data_col135[103] <= data_col135[102];
   data_col135[104] <= data_col135[103];
   data_col135[105] <= data_col135[104];
   data_col135[106] <= data_col135[105];
   data_col135[107] <= data_col135[106];
   data_col135[108] <= data_col135[107];
   data_col135[109] <= data_col135[108];
   data_col135[110] <= data_col135[109];
   data_col135[111] <= data_col135[110];
   data_col135[112] <= data_col135[111];
   data_col135[113] <= data_col135[112];
   data_col135[114] <= data_col135[113];
   data_col135[115] <= data_col135[114];
   data_col135[116] <= data_col135[115];
   data_col135[117] <= data_col135[116];
   data_col135[118] <= data_col135[117];
   data_col135[119] <= data_col135[118];
   data_col135[120] <= data_col135[119];
   data_col135[121] <= data_col135[120];
   data_col135[122] <= data_col135[121];
   data_col135[123] <= data_col135[122];
   data_col135[124] <= data_col135[123];
   data_col135[125] <= data_col135[124];
   data_col135[126] <= data_col135[125];
   data_col135[127] <= data_col135[126];
   data_col135[128] <= data_col135[127];
   data_col135[129] <= data_col135[128];
   data_col135[130] <= data_col135[129];
   data_col135[131] <= data_col135[130];
   data_col135[132] <= data_col135[131];
   data_col135[133] <= data_col135[132];
   data_col135[134] <= data_col135[133];
   data_col135[135] <= data_col135[134];

   data_col136[1] <= data[29];
   data_col136[2] <= data_col136[1];
   data_col136[3] <= data_col136[2];
   data_col136[4] <= data_col136[3];
   data_col136[5] <= data_col136[4];
   data_col136[6] <= data_col136[5];
   data_col136[7] <= data_col136[6];
   data_col136[8] <= data_col136[7];
   data_col136[9] <= data_col136[8];
   data_col136[10] <= data_col136[9];
   data_col136[11] <= data_col136[10];
   data_col136[12] <= data_col136[11];
   data_col136[13] <= data_col136[12];
   data_col136[14] <= data_col136[13];
   data_col136[15] <= data_col136[14];
   data_col136[16] <= data_col136[15];
   data_col136[17] <= data_col136[16];
   data_col136[18] <= data_col136[17];
   data_col136[19] <= data_col136[18];
   data_col136[20] <= data_col136[19];
   data_col136[21] <= data_col136[20];
   data_col136[22] <= data_col136[21];
   data_col136[23] <= data_col136[22];
   data_col136[24] <= data_col136[23];
   data_col136[25] <= data_col136[24];
   data_col136[26] <= data_col136[25];
   data_col136[27] <= data_col136[26];
   data_col136[28] <= data_col136[27];
   data_col136[29] <= data_col136[28];
   data_col136[30] <= data_col136[29];
   data_col136[31] <= data_col136[30];
   data_col136[32] <= data_col136[31];
   data_col136[33] <= data_col136[32];
   data_col136[34] <= data_col136[33];
   data_col136[35] <= data_col136[34];
   data_col136[36] <= data_col136[35];
   data_col136[37] <= data_col136[36];
   data_col136[38] <= data_col136[37];
   data_col136[39] <= data_col136[38];
   data_col136[40] <= data_col136[39];
   data_col136[41] <= data_col136[40];
   data_col136[42] <= data_col136[41];
   data_col136[43] <= data_col136[42];
   data_col136[44] <= data_col136[43];
   data_col136[45] <= data_col136[44];
   data_col136[46] <= data_col136[45];
   data_col136[47] <= data_col136[46];
   data_col136[48] <= data_col136[47];
   data_col136[49] <= data_col136[48];
   data_col136[50] <= data_col136[49];
   data_col136[51] <= data_col136[50];
   data_col136[52] <= data_col136[51];
   data_col136[53] <= data_col136[52];
   data_col136[54] <= data_col136[53];
   data_col136[55] <= data_col136[54];
   data_col136[56] <= data_col136[55];
   data_col136[57] <= data_col136[56];
   data_col136[58] <= data_col136[57];
   data_col136[59] <= data_col136[58];
   data_col136[60] <= data_col136[59];
   data_col136[61] <= data_col136[60];
   data_col136[62] <= data_col136[61];
   data_col136[63] <= data_col136[62];
   data_col136[64] <= data_col136[63];
   data_col136[65] <= data_col136[64];
   data_col136[66] <= data_col136[65];
   data_col136[67] <= data_col136[66];
   data_col136[68] <= data_col136[67];
   data_col136[69] <= data_col136[68];
   data_col136[70] <= data_col136[69];
   data_col136[71] <= data_col136[70];
   data_col136[72] <= data_col136[71];
   data_col136[73] <= data_col136[72];
   data_col136[74] <= data_col136[73];
   data_col136[75] <= data_col136[74];
   data_col136[76] <= data_col136[75];
   data_col136[77] <= data_col136[76];
   data_col136[78] <= data_col136[77];
   data_col136[79] <= data_col136[78];
   data_col136[80] <= data_col136[79];
   data_col136[81] <= data_col136[80];
   data_col136[82] <= data_col136[81];
   data_col136[83] <= data_col136[82];
   data_col136[84] <= data_col136[83];
   data_col136[85] <= data_col136[84];
   data_col136[86] <= data_col136[85];
   data_col136[87] <= data_col136[86];
   data_col136[88] <= data_col136[87];
   data_col136[89] <= data_col136[88];
   data_col136[90] <= data_col136[89];
   data_col136[91] <= data_col136[90];
   data_col136[92] <= data_col136[91];
   data_col136[93] <= data_col136[92];
   data_col136[94] <= data_col136[93];
   data_col136[95] <= data_col136[94];
   data_col136[96] <= data_col136[95];
   data_col136[97] <= data_col136[96];
   data_col136[98] <= data_col136[97];
   data_col136[99] <= data_col136[98];
   data_col136[100] <= data_col136[99];
   data_col136[101] <= data_col136[100];
   data_col136[102] <= data_col136[101];
   data_col136[103] <= data_col136[102];
   data_col136[104] <= data_col136[103];
   data_col136[105] <= data_col136[104];
   data_col136[106] <= data_col136[105];
   data_col136[107] <= data_col136[106];
   data_col136[108] <= data_col136[107];
   data_col136[109] <= data_col136[108];
   data_col136[110] <= data_col136[109];
   data_col136[111] <= data_col136[110];
   data_col136[112] <= data_col136[111];
   data_col136[113] <= data_col136[112];
   data_col136[114] <= data_col136[113];
   data_col136[115] <= data_col136[114];
   data_col136[116] <= data_col136[115];
   data_col136[117] <= data_col136[116];
   data_col136[118] <= data_col136[117];
   data_col136[119] <= data_col136[118];
   data_col136[120] <= data_col136[119];
   data_col136[121] <= data_col136[120];
   data_col136[122] <= data_col136[121];
   data_col136[123] <= data_col136[122];
   data_col136[124] <= data_col136[123];
   data_col136[125] <= data_col136[124];
   data_col136[126] <= data_col136[125];
   data_col136[127] <= data_col136[126];
   data_col136[128] <= data_col136[127];
   data_col136[129] <= data_col136[128];
   data_col136[130] <= data_col136[129];
   data_col136[131] <= data_col136[130];
   data_col136[132] <= data_col136[131];
   data_col136[133] <= data_col136[132];
   data_col136[134] <= data_col136[133];
   data_col136[135] <= data_col136[134];
   data_col136[136] <= data_col136[135];

   data_col137[1] <= data[28];
   data_col137[2] <= data_col137[1];
   data_col137[3] <= data_col137[2];
   data_col137[4] <= data_col137[3];
   data_col137[5] <= data_col137[4];
   data_col137[6] <= data_col137[5];
   data_col137[7] <= data_col137[6];
   data_col137[8] <= data_col137[7];
   data_col137[9] <= data_col137[8];
   data_col137[10] <= data_col137[9];
   data_col137[11] <= data_col137[10];
   data_col137[12] <= data_col137[11];
   data_col137[13] <= data_col137[12];
   data_col137[14] <= data_col137[13];
   data_col137[15] <= data_col137[14];
   data_col137[16] <= data_col137[15];
   data_col137[17] <= data_col137[16];
   data_col137[18] <= data_col137[17];
   data_col137[19] <= data_col137[18];
   data_col137[20] <= data_col137[19];
   data_col137[21] <= data_col137[20];
   data_col137[22] <= data_col137[21];
   data_col137[23] <= data_col137[22];
   data_col137[24] <= data_col137[23];
   data_col137[25] <= data_col137[24];
   data_col137[26] <= data_col137[25];
   data_col137[27] <= data_col137[26];
   data_col137[28] <= data_col137[27];
   data_col137[29] <= data_col137[28];
   data_col137[30] <= data_col137[29];
   data_col137[31] <= data_col137[30];
   data_col137[32] <= data_col137[31];
   data_col137[33] <= data_col137[32];
   data_col137[34] <= data_col137[33];
   data_col137[35] <= data_col137[34];
   data_col137[36] <= data_col137[35];
   data_col137[37] <= data_col137[36];
   data_col137[38] <= data_col137[37];
   data_col137[39] <= data_col137[38];
   data_col137[40] <= data_col137[39];
   data_col137[41] <= data_col137[40];
   data_col137[42] <= data_col137[41];
   data_col137[43] <= data_col137[42];
   data_col137[44] <= data_col137[43];
   data_col137[45] <= data_col137[44];
   data_col137[46] <= data_col137[45];
   data_col137[47] <= data_col137[46];
   data_col137[48] <= data_col137[47];
   data_col137[49] <= data_col137[48];
   data_col137[50] <= data_col137[49];
   data_col137[51] <= data_col137[50];
   data_col137[52] <= data_col137[51];
   data_col137[53] <= data_col137[52];
   data_col137[54] <= data_col137[53];
   data_col137[55] <= data_col137[54];
   data_col137[56] <= data_col137[55];
   data_col137[57] <= data_col137[56];
   data_col137[58] <= data_col137[57];
   data_col137[59] <= data_col137[58];
   data_col137[60] <= data_col137[59];
   data_col137[61] <= data_col137[60];
   data_col137[62] <= data_col137[61];
   data_col137[63] <= data_col137[62];
   data_col137[64] <= data_col137[63];
   data_col137[65] <= data_col137[64];
   data_col137[66] <= data_col137[65];
   data_col137[67] <= data_col137[66];
   data_col137[68] <= data_col137[67];
   data_col137[69] <= data_col137[68];
   data_col137[70] <= data_col137[69];
   data_col137[71] <= data_col137[70];
   data_col137[72] <= data_col137[71];
   data_col137[73] <= data_col137[72];
   data_col137[74] <= data_col137[73];
   data_col137[75] <= data_col137[74];
   data_col137[76] <= data_col137[75];
   data_col137[77] <= data_col137[76];
   data_col137[78] <= data_col137[77];
   data_col137[79] <= data_col137[78];
   data_col137[80] <= data_col137[79];
   data_col137[81] <= data_col137[80];
   data_col137[82] <= data_col137[81];
   data_col137[83] <= data_col137[82];
   data_col137[84] <= data_col137[83];
   data_col137[85] <= data_col137[84];
   data_col137[86] <= data_col137[85];
   data_col137[87] <= data_col137[86];
   data_col137[88] <= data_col137[87];
   data_col137[89] <= data_col137[88];
   data_col137[90] <= data_col137[89];
   data_col137[91] <= data_col137[90];
   data_col137[92] <= data_col137[91];
   data_col137[93] <= data_col137[92];
   data_col137[94] <= data_col137[93];
   data_col137[95] <= data_col137[94];
   data_col137[96] <= data_col137[95];
   data_col137[97] <= data_col137[96];
   data_col137[98] <= data_col137[97];
   data_col137[99] <= data_col137[98];
   data_col137[100] <= data_col137[99];
   data_col137[101] <= data_col137[100];
   data_col137[102] <= data_col137[101];
   data_col137[103] <= data_col137[102];
   data_col137[104] <= data_col137[103];
   data_col137[105] <= data_col137[104];
   data_col137[106] <= data_col137[105];
   data_col137[107] <= data_col137[106];
   data_col137[108] <= data_col137[107];
   data_col137[109] <= data_col137[108];
   data_col137[110] <= data_col137[109];
   data_col137[111] <= data_col137[110];
   data_col137[112] <= data_col137[111];
   data_col137[113] <= data_col137[112];
   data_col137[114] <= data_col137[113];
   data_col137[115] <= data_col137[114];
   data_col137[116] <= data_col137[115];
   data_col137[117] <= data_col137[116];
   data_col137[118] <= data_col137[117];
   data_col137[119] <= data_col137[118];
   data_col137[120] <= data_col137[119];
   data_col137[121] <= data_col137[120];
   data_col137[122] <= data_col137[121];
   data_col137[123] <= data_col137[122];
   data_col137[124] <= data_col137[123];
   data_col137[125] <= data_col137[124];
   data_col137[126] <= data_col137[125];
   data_col137[127] <= data_col137[126];
   data_col137[128] <= data_col137[127];
   data_col137[129] <= data_col137[128];
   data_col137[130] <= data_col137[129];
   data_col137[131] <= data_col137[130];
   data_col137[132] <= data_col137[131];
   data_col137[133] <= data_col137[132];
   data_col137[134] <= data_col137[133];
   data_col137[135] <= data_col137[134];
   data_col137[136] <= data_col137[135];
   data_col137[137] <= data_col137[136];

   data_col138[1] <= data[27];
   data_col138[2] <= data_col138[1];
   data_col138[3] <= data_col138[2];
   data_col138[4] <= data_col138[3];
   data_col138[5] <= data_col138[4];
   data_col138[6] <= data_col138[5];
   data_col138[7] <= data_col138[6];
   data_col138[8] <= data_col138[7];
   data_col138[9] <= data_col138[8];
   data_col138[10] <= data_col138[9];
   data_col138[11] <= data_col138[10];
   data_col138[12] <= data_col138[11];
   data_col138[13] <= data_col138[12];
   data_col138[14] <= data_col138[13];
   data_col138[15] <= data_col138[14];
   data_col138[16] <= data_col138[15];
   data_col138[17] <= data_col138[16];
   data_col138[18] <= data_col138[17];
   data_col138[19] <= data_col138[18];
   data_col138[20] <= data_col138[19];
   data_col138[21] <= data_col138[20];
   data_col138[22] <= data_col138[21];
   data_col138[23] <= data_col138[22];
   data_col138[24] <= data_col138[23];
   data_col138[25] <= data_col138[24];
   data_col138[26] <= data_col138[25];
   data_col138[27] <= data_col138[26];
   data_col138[28] <= data_col138[27];
   data_col138[29] <= data_col138[28];
   data_col138[30] <= data_col138[29];
   data_col138[31] <= data_col138[30];
   data_col138[32] <= data_col138[31];
   data_col138[33] <= data_col138[32];
   data_col138[34] <= data_col138[33];
   data_col138[35] <= data_col138[34];
   data_col138[36] <= data_col138[35];
   data_col138[37] <= data_col138[36];
   data_col138[38] <= data_col138[37];
   data_col138[39] <= data_col138[38];
   data_col138[40] <= data_col138[39];
   data_col138[41] <= data_col138[40];
   data_col138[42] <= data_col138[41];
   data_col138[43] <= data_col138[42];
   data_col138[44] <= data_col138[43];
   data_col138[45] <= data_col138[44];
   data_col138[46] <= data_col138[45];
   data_col138[47] <= data_col138[46];
   data_col138[48] <= data_col138[47];
   data_col138[49] <= data_col138[48];
   data_col138[50] <= data_col138[49];
   data_col138[51] <= data_col138[50];
   data_col138[52] <= data_col138[51];
   data_col138[53] <= data_col138[52];
   data_col138[54] <= data_col138[53];
   data_col138[55] <= data_col138[54];
   data_col138[56] <= data_col138[55];
   data_col138[57] <= data_col138[56];
   data_col138[58] <= data_col138[57];
   data_col138[59] <= data_col138[58];
   data_col138[60] <= data_col138[59];
   data_col138[61] <= data_col138[60];
   data_col138[62] <= data_col138[61];
   data_col138[63] <= data_col138[62];
   data_col138[64] <= data_col138[63];
   data_col138[65] <= data_col138[64];
   data_col138[66] <= data_col138[65];
   data_col138[67] <= data_col138[66];
   data_col138[68] <= data_col138[67];
   data_col138[69] <= data_col138[68];
   data_col138[70] <= data_col138[69];
   data_col138[71] <= data_col138[70];
   data_col138[72] <= data_col138[71];
   data_col138[73] <= data_col138[72];
   data_col138[74] <= data_col138[73];
   data_col138[75] <= data_col138[74];
   data_col138[76] <= data_col138[75];
   data_col138[77] <= data_col138[76];
   data_col138[78] <= data_col138[77];
   data_col138[79] <= data_col138[78];
   data_col138[80] <= data_col138[79];
   data_col138[81] <= data_col138[80];
   data_col138[82] <= data_col138[81];
   data_col138[83] <= data_col138[82];
   data_col138[84] <= data_col138[83];
   data_col138[85] <= data_col138[84];
   data_col138[86] <= data_col138[85];
   data_col138[87] <= data_col138[86];
   data_col138[88] <= data_col138[87];
   data_col138[89] <= data_col138[88];
   data_col138[90] <= data_col138[89];
   data_col138[91] <= data_col138[90];
   data_col138[92] <= data_col138[91];
   data_col138[93] <= data_col138[92];
   data_col138[94] <= data_col138[93];
   data_col138[95] <= data_col138[94];
   data_col138[96] <= data_col138[95];
   data_col138[97] <= data_col138[96];
   data_col138[98] <= data_col138[97];
   data_col138[99] <= data_col138[98];
   data_col138[100] <= data_col138[99];
   data_col138[101] <= data_col138[100];
   data_col138[102] <= data_col138[101];
   data_col138[103] <= data_col138[102];
   data_col138[104] <= data_col138[103];
   data_col138[105] <= data_col138[104];
   data_col138[106] <= data_col138[105];
   data_col138[107] <= data_col138[106];
   data_col138[108] <= data_col138[107];
   data_col138[109] <= data_col138[108];
   data_col138[110] <= data_col138[109];
   data_col138[111] <= data_col138[110];
   data_col138[112] <= data_col138[111];
   data_col138[113] <= data_col138[112];
   data_col138[114] <= data_col138[113];
   data_col138[115] <= data_col138[114];
   data_col138[116] <= data_col138[115];
   data_col138[117] <= data_col138[116];
   data_col138[118] <= data_col138[117];
   data_col138[119] <= data_col138[118];
   data_col138[120] <= data_col138[119];
   data_col138[121] <= data_col138[120];
   data_col138[122] <= data_col138[121];
   data_col138[123] <= data_col138[122];
   data_col138[124] <= data_col138[123];
   data_col138[125] <= data_col138[124];
   data_col138[126] <= data_col138[125];
   data_col138[127] <= data_col138[126];
   data_col138[128] <= data_col138[127];
   data_col138[129] <= data_col138[128];
   data_col138[130] <= data_col138[129];
   data_col138[131] <= data_col138[130];
   data_col138[132] <= data_col138[131];
   data_col138[133] <= data_col138[132];
   data_col138[134] <= data_col138[133];
   data_col138[135] <= data_col138[134];
   data_col138[136] <= data_col138[135];
   data_col138[137] <= data_col138[136];
   data_col138[138] <= data_col138[137];

   data_col139[1] <= data[26];
   data_col139[2] <= data_col139[1];
   data_col139[3] <= data_col139[2];
   data_col139[4] <= data_col139[3];
   data_col139[5] <= data_col139[4];
   data_col139[6] <= data_col139[5];
   data_col139[7] <= data_col139[6];
   data_col139[8] <= data_col139[7];
   data_col139[9] <= data_col139[8];
   data_col139[10] <= data_col139[9];
   data_col139[11] <= data_col139[10];
   data_col139[12] <= data_col139[11];
   data_col139[13] <= data_col139[12];
   data_col139[14] <= data_col139[13];
   data_col139[15] <= data_col139[14];
   data_col139[16] <= data_col139[15];
   data_col139[17] <= data_col139[16];
   data_col139[18] <= data_col139[17];
   data_col139[19] <= data_col139[18];
   data_col139[20] <= data_col139[19];
   data_col139[21] <= data_col139[20];
   data_col139[22] <= data_col139[21];
   data_col139[23] <= data_col139[22];
   data_col139[24] <= data_col139[23];
   data_col139[25] <= data_col139[24];
   data_col139[26] <= data_col139[25];
   data_col139[27] <= data_col139[26];
   data_col139[28] <= data_col139[27];
   data_col139[29] <= data_col139[28];
   data_col139[30] <= data_col139[29];
   data_col139[31] <= data_col139[30];
   data_col139[32] <= data_col139[31];
   data_col139[33] <= data_col139[32];
   data_col139[34] <= data_col139[33];
   data_col139[35] <= data_col139[34];
   data_col139[36] <= data_col139[35];
   data_col139[37] <= data_col139[36];
   data_col139[38] <= data_col139[37];
   data_col139[39] <= data_col139[38];
   data_col139[40] <= data_col139[39];
   data_col139[41] <= data_col139[40];
   data_col139[42] <= data_col139[41];
   data_col139[43] <= data_col139[42];
   data_col139[44] <= data_col139[43];
   data_col139[45] <= data_col139[44];
   data_col139[46] <= data_col139[45];
   data_col139[47] <= data_col139[46];
   data_col139[48] <= data_col139[47];
   data_col139[49] <= data_col139[48];
   data_col139[50] <= data_col139[49];
   data_col139[51] <= data_col139[50];
   data_col139[52] <= data_col139[51];
   data_col139[53] <= data_col139[52];
   data_col139[54] <= data_col139[53];
   data_col139[55] <= data_col139[54];
   data_col139[56] <= data_col139[55];
   data_col139[57] <= data_col139[56];
   data_col139[58] <= data_col139[57];
   data_col139[59] <= data_col139[58];
   data_col139[60] <= data_col139[59];
   data_col139[61] <= data_col139[60];
   data_col139[62] <= data_col139[61];
   data_col139[63] <= data_col139[62];
   data_col139[64] <= data_col139[63];
   data_col139[65] <= data_col139[64];
   data_col139[66] <= data_col139[65];
   data_col139[67] <= data_col139[66];
   data_col139[68] <= data_col139[67];
   data_col139[69] <= data_col139[68];
   data_col139[70] <= data_col139[69];
   data_col139[71] <= data_col139[70];
   data_col139[72] <= data_col139[71];
   data_col139[73] <= data_col139[72];
   data_col139[74] <= data_col139[73];
   data_col139[75] <= data_col139[74];
   data_col139[76] <= data_col139[75];
   data_col139[77] <= data_col139[76];
   data_col139[78] <= data_col139[77];
   data_col139[79] <= data_col139[78];
   data_col139[80] <= data_col139[79];
   data_col139[81] <= data_col139[80];
   data_col139[82] <= data_col139[81];
   data_col139[83] <= data_col139[82];
   data_col139[84] <= data_col139[83];
   data_col139[85] <= data_col139[84];
   data_col139[86] <= data_col139[85];
   data_col139[87] <= data_col139[86];
   data_col139[88] <= data_col139[87];
   data_col139[89] <= data_col139[88];
   data_col139[90] <= data_col139[89];
   data_col139[91] <= data_col139[90];
   data_col139[92] <= data_col139[91];
   data_col139[93] <= data_col139[92];
   data_col139[94] <= data_col139[93];
   data_col139[95] <= data_col139[94];
   data_col139[96] <= data_col139[95];
   data_col139[97] <= data_col139[96];
   data_col139[98] <= data_col139[97];
   data_col139[99] <= data_col139[98];
   data_col139[100] <= data_col139[99];
   data_col139[101] <= data_col139[100];
   data_col139[102] <= data_col139[101];
   data_col139[103] <= data_col139[102];
   data_col139[104] <= data_col139[103];
   data_col139[105] <= data_col139[104];
   data_col139[106] <= data_col139[105];
   data_col139[107] <= data_col139[106];
   data_col139[108] <= data_col139[107];
   data_col139[109] <= data_col139[108];
   data_col139[110] <= data_col139[109];
   data_col139[111] <= data_col139[110];
   data_col139[112] <= data_col139[111];
   data_col139[113] <= data_col139[112];
   data_col139[114] <= data_col139[113];
   data_col139[115] <= data_col139[114];
   data_col139[116] <= data_col139[115];
   data_col139[117] <= data_col139[116];
   data_col139[118] <= data_col139[117];
   data_col139[119] <= data_col139[118];
   data_col139[120] <= data_col139[119];
   data_col139[121] <= data_col139[120];
   data_col139[122] <= data_col139[121];
   data_col139[123] <= data_col139[122];
   data_col139[124] <= data_col139[123];
   data_col139[125] <= data_col139[124];
   data_col139[126] <= data_col139[125];
   data_col139[127] <= data_col139[126];
   data_col139[128] <= data_col139[127];
   data_col139[129] <= data_col139[128];
   data_col139[130] <= data_col139[129];
   data_col139[131] <= data_col139[130];
   data_col139[132] <= data_col139[131];
   data_col139[133] <= data_col139[132];
   data_col139[134] <= data_col139[133];
   data_col139[135] <= data_col139[134];
   data_col139[136] <= data_col139[135];
   data_col139[137] <= data_col139[136];
   data_col139[138] <= data_col139[137];
   data_col139[139] <= data_col139[138];

   data_col140[1] <= data[25];
   data_col140[2] <= data_col140[1];
   data_col140[3] <= data_col140[2];
   data_col140[4] <= data_col140[3];
   data_col140[5] <= data_col140[4];
   data_col140[6] <= data_col140[5];
   data_col140[7] <= data_col140[6];
   data_col140[8] <= data_col140[7];
   data_col140[9] <= data_col140[8];
   data_col140[10] <= data_col140[9];
   data_col140[11] <= data_col140[10];
   data_col140[12] <= data_col140[11];
   data_col140[13] <= data_col140[12];
   data_col140[14] <= data_col140[13];
   data_col140[15] <= data_col140[14];
   data_col140[16] <= data_col140[15];
   data_col140[17] <= data_col140[16];
   data_col140[18] <= data_col140[17];
   data_col140[19] <= data_col140[18];
   data_col140[20] <= data_col140[19];
   data_col140[21] <= data_col140[20];
   data_col140[22] <= data_col140[21];
   data_col140[23] <= data_col140[22];
   data_col140[24] <= data_col140[23];
   data_col140[25] <= data_col140[24];
   data_col140[26] <= data_col140[25];
   data_col140[27] <= data_col140[26];
   data_col140[28] <= data_col140[27];
   data_col140[29] <= data_col140[28];
   data_col140[30] <= data_col140[29];
   data_col140[31] <= data_col140[30];
   data_col140[32] <= data_col140[31];
   data_col140[33] <= data_col140[32];
   data_col140[34] <= data_col140[33];
   data_col140[35] <= data_col140[34];
   data_col140[36] <= data_col140[35];
   data_col140[37] <= data_col140[36];
   data_col140[38] <= data_col140[37];
   data_col140[39] <= data_col140[38];
   data_col140[40] <= data_col140[39];
   data_col140[41] <= data_col140[40];
   data_col140[42] <= data_col140[41];
   data_col140[43] <= data_col140[42];
   data_col140[44] <= data_col140[43];
   data_col140[45] <= data_col140[44];
   data_col140[46] <= data_col140[45];
   data_col140[47] <= data_col140[46];
   data_col140[48] <= data_col140[47];
   data_col140[49] <= data_col140[48];
   data_col140[50] <= data_col140[49];
   data_col140[51] <= data_col140[50];
   data_col140[52] <= data_col140[51];
   data_col140[53] <= data_col140[52];
   data_col140[54] <= data_col140[53];
   data_col140[55] <= data_col140[54];
   data_col140[56] <= data_col140[55];
   data_col140[57] <= data_col140[56];
   data_col140[58] <= data_col140[57];
   data_col140[59] <= data_col140[58];
   data_col140[60] <= data_col140[59];
   data_col140[61] <= data_col140[60];
   data_col140[62] <= data_col140[61];
   data_col140[63] <= data_col140[62];
   data_col140[64] <= data_col140[63];
   data_col140[65] <= data_col140[64];
   data_col140[66] <= data_col140[65];
   data_col140[67] <= data_col140[66];
   data_col140[68] <= data_col140[67];
   data_col140[69] <= data_col140[68];
   data_col140[70] <= data_col140[69];
   data_col140[71] <= data_col140[70];
   data_col140[72] <= data_col140[71];
   data_col140[73] <= data_col140[72];
   data_col140[74] <= data_col140[73];
   data_col140[75] <= data_col140[74];
   data_col140[76] <= data_col140[75];
   data_col140[77] <= data_col140[76];
   data_col140[78] <= data_col140[77];
   data_col140[79] <= data_col140[78];
   data_col140[80] <= data_col140[79];
   data_col140[81] <= data_col140[80];
   data_col140[82] <= data_col140[81];
   data_col140[83] <= data_col140[82];
   data_col140[84] <= data_col140[83];
   data_col140[85] <= data_col140[84];
   data_col140[86] <= data_col140[85];
   data_col140[87] <= data_col140[86];
   data_col140[88] <= data_col140[87];
   data_col140[89] <= data_col140[88];
   data_col140[90] <= data_col140[89];
   data_col140[91] <= data_col140[90];
   data_col140[92] <= data_col140[91];
   data_col140[93] <= data_col140[92];
   data_col140[94] <= data_col140[93];
   data_col140[95] <= data_col140[94];
   data_col140[96] <= data_col140[95];
   data_col140[97] <= data_col140[96];
   data_col140[98] <= data_col140[97];
   data_col140[99] <= data_col140[98];
   data_col140[100] <= data_col140[99];
   data_col140[101] <= data_col140[100];
   data_col140[102] <= data_col140[101];
   data_col140[103] <= data_col140[102];
   data_col140[104] <= data_col140[103];
   data_col140[105] <= data_col140[104];
   data_col140[106] <= data_col140[105];
   data_col140[107] <= data_col140[106];
   data_col140[108] <= data_col140[107];
   data_col140[109] <= data_col140[108];
   data_col140[110] <= data_col140[109];
   data_col140[111] <= data_col140[110];
   data_col140[112] <= data_col140[111];
   data_col140[113] <= data_col140[112];
   data_col140[114] <= data_col140[113];
   data_col140[115] <= data_col140[114];
   data_col140[116] <= data_col140[115];
   data_col140[117] <= data_col140[116];
   data_col140[118] <= data_col140[117];
   data_col140[119] <= data_col140[118];
   data_col140[120] <= data_col140[119];
   data_col140[121] <= data_col140[120];
   data_col140[122] <= data_col140[121];
   data_col140[123] <= data_col140[122];
   data_col140[124] <= data_col140[123];
   data_col140[125] <= data_col140[124];
   data_col140[126] <= data_col140[125];
   data_col140[127] <= data_col140[126];
   data_col140[128] <= data_col140[127];
   data_col140[129] <= data_col140[128];
   data_col140[130] <= data_col140[129];
   data_col140[131] <= data_col140[130];
   data_col140[132] <= data_col140[131];
   data_col140[133] <= data_col140[132];
   data_col140[134] <= data_col140[133];
   data_col140[135] <= data_col140[134];
   data_col140[136] <= data_col140[135];
   data_col140[137] <= data_col140[136];
   data_col140[138] <= data_col140[137];
   data_col140[139] <= data_col140[138];
   data_col140[140] <= data_col140[139];

   data_col141[1] <= data[24];
   data_col141[2] <= data_col141[1];
   data_col141[3] <= data_col141[2];
   data_col141[4] <= data_col141[3];
   data_col141[5] <= data_col141[4];
   data_col141[6] <= data_col141[5];
   data_col141[7] <= data_col141[6];
   data_col141[8] <= data_col141[7];
   data_col141[9] <= data_col141[8];
   data_col141[10] <= data_col141[9];
   data_col141[11] <= data_col141[10];
   data_col141[12] <= data_col141[11];
   data_col141[13] <= data_col141[12];
   data_col141[14] <= data_col141[13];
   data_col141[15] <= data_col141[14];
   data_col141[16] <= data_col141[15];
   data_col141[17] <= data_col141[16];
   data_col141[18] <= data_col141[17];
   data_col141[19] <= data_col141[18];
   data_col141[20] <= data_col141[19];
   data_col141[21] <= data_col141[20];
   data_col141[22] <= data_col141[21];
   data_col141[23] <= data_col141[22];
   data_col141[24] <= data_col141[23];
   data_col141[25] <= data_col141[24];
   data_col141[26] <= data_col141[25];
   data_col141[27] <= data_col141[26];
   data_col141[28] <= data_col141[27];
   data_col141[29] <= data_col141[28];
   data_col141[30] <= data_col141[29];
   data_col141[31] <= data_col141[30];
   data_col141[32] <= data_col141[31];
   data_col141[33] <= data_col141[32];
   data_col141[34] <= data_col141[33];
   data_col141[35] <= data_col141[34];
   data_col141[36] <= data_col141[35];
   data_col141[37] <= data_col141[36];
   data_col141[38] <= data_col141[37];
   data_col141[39] <= data_col141[38];
   data_col141[40] <= data_col141[39];
   data_col141[41] <= data_col141[40];
   data_col141[42] <= data_col141[41];
   data_col141[43] <= data_col141[42];
   data_col141[44] <= data_col141[43];
   data_col141[45] <= data_col141[44];
   data_col141[46] <= data_col141[45];
   data_col141[47] <= data_col141[46];
   data_col141[48] <= data_col141[47];
   data_col141[49] <= data_col141[48];
   data_col141[50] <= data_col141[49];
   data_col141[51] <= data_col141[50];
   data_col141[52] <= data_col141[51];
   data_col141[53] <= data_col141[52];
   data_col141[54] <= data_col141[53];
   data_col141[55] <= data_col141[54];
   data_col141[56] <= data_col141[55];
   data_col141[57] <= data_col141[56];
   data_col141[58] <= data_col141[57];
   data_col141[59] <= data_col141[58];
   data_col141[60] <= data_col141[59];
   data_col141[61] <= data_col141[60];
   data_col141[62] <= data_col141[61];
   data_col141[63] <= data_col141[62];
   data_col141[64] <= data_col141[63];
   data_col141[65] <= data_col141[64];
   data_col141[66] <= data_col141[65];
   data_col141[67] <= data_col141[66];
   data_col141[68] <= data_col141[67];
   data_col141[69] <= data_col141[68];
   data_col141[70] <= data_col141[69];
   data_col141[71] <= data_col141[70];
   data_col141[72] <= data_col141[71];
   data_col141[73] <= data_col141[72];
   data_col141[74] <= data_col141[73];
   data_col141[75] <= data_col141[74];
   data_col141[76] <= data_col141[75];
   data_col141[77] <= data_col141[76];
   data_col141[78] <= data_col141[77];
   data_col141[79] <= data_col141[78];
   data_col141[80] <= data_col141[79];
   data_col141[81] <= data_col141[80];
   data_col141[82] <= data_col141[81];
   data_col141[83] <= data_col141[82];
   data_col141[84] <= data_col141[83];
   data_col141[85] <= data_col141[84];
   data_col141[86] <= data_col141[85];
   data_col141[87] <= data_col141[86];
   data_col141[88] <= data_col141[87];
   data_col141[89] <= data_col141[88];
   data_col141[90] <= data_col141[89];
   data_col141[91] <= data_col141[90];
   data_col141[92] <= data_col141[91];
   data_col141[93] <= data_col141[92];
   data_col141[94] <= data_col141[93];
   data_col141[95] <= data_col141[94];
   data_col141[96] <= data_col141[95];
   data_col141[97] <= data_col141[96];
   data_col141[98] <= data_col141[97];
   data_col141[99] <= data_col141[98];
   data_col141[100] <= data_col141[99];
   data_col141[101] <= data_col141[100];
   data_col141[102] <= data_col141[101];
   data_col141[103] <= data_col141[102];
   data_col141[104] <= data_col141[103];
   data_col141[105] <= data_col141[104];
   data_col141[106] <= data_col141[105];
   data_col141[107] <= data_col141[106];
   data_col141[108] <= data_col141[107];
   data_col141[109] <= data_col141[108];
   data_col141[110] <= data_col141[109];
   data_col141[111] <= data_col141[110];
   data_col141[112] <= data_col141[111];
   data_col141[113] <= data_col141[112];
   data_col141[114] <= data_col141[113];
   data_col141[115] <= data_col141[114];
   data_col141[116] <= data_col141[115];
   data_col141[117] <= data_col141[116];
   data_col141[118] <= data_col141[117];
   data_col141[119] <= data_col141[118];
   data_col141[120] <= data_col141[119];
   data_col141[121] <= data_col141[120];
   data_col141[122] <= data_col141[121];
   data_col141[123] <= data_col141[122];
   data_col141[124] <= data_col141[123];
   data_col141[125] <= data_col141[124];
   data_col141[126] <= data_col141[125];
   data_col141[127] <= data_col141[126];
   data_col141[128] <= data_col141[127];
   data_col141[129] <= data_col141[128];
   data_col141[130] <= data_col141[129];
   data_col141[131] <= data_col141[130];
   data_col141[132] <= data_col141[131];
   data_col141[133] <= data_col141[132];
   data_col141[134] <= data_col141[133];
   data_col141[135] <= data_col141[134];
   data_col141[136] <= data_col141[135];
   data_col141[137] <= data_col141[136];
   data_col141[138] <= data_col141[137];
   data_col141[139] <= data_col141[138];
   data_col141[140] <= data_col141[139];
   data_col141[141] <= data_col141[140];

   data_col142[1] <= data[23];
   data_col142[2] <= data_col142[1];
   data_col142[3] <= data_col142[2];
   data_col142[4] <= data_col142[3];
   data_col142[5] <= data_col142[4];
   data_col142[6] <= data_col142[5];
   data_col142[7] <= data_col142[6];
   data_col142[8] <= data_col142[7];
   data_col142[9] <= data_col142[8];
   data_col142[10] <= data_col142[9];
   data_col142[11] <= data_col142[10];
   data_col142[12] <= data_col142[11];
   data_col142[13] <= data_col142[12];
   data_col142[14] <= data_col142[13];
   data_col142[15] <= data_col142[14];
   data_col142[16] <= data_col142[15];
   data_col142[17] <= data_col142[16];
   data_col142[18] <= data_col142[17];
   data_col142[19] <= data_col142[18];
   data_col142[20] <= data_col142[19];
   data_col142[21] <= data_col142[20];
   data_col142[22] <= data_col142[21];
   data_col142[23] <= data_col142[22];
   data_col142[24] <= data_col142[23];
   data_col142[25] <= data_col142[24];
   data_col142[26] <= data_col142[25];
   data_col142[27] <= data_col142[26];
   data_col142[28] <= data_col142[27];
   data_col142[29] <= data_col142[28];
   data_col142[30] <= data_col142[29];
   data_col142[31] <= data_col142[30];
   data_col142[32] <= data_col142[31];
   data_col142[33] <= data_col142[32];
   data_col142[34] <= data_col142[33];
   data_col142[35] <= data_col142[34];
   data_col142[36] <= data_col142[35];
   data_col142[37] <= data_col142[36];
   data_col142[38] <= data_col142[37];
   data_col142[39] <= data_col142[38];
   data_col142[40] <= data_col142[39];
   data_col142[41] <= data_col142[40];
   data_col142[42] <= data_col142[41];
   data_col142[43] <= data_col142[42];
   data_col142[44] <= data_col142[43];
   data_col142[45] <= data_col142[44];
   data_col142[46] <= data_col142[45];
   data_col142[47] <= data_col142[46];
   data_col142[48] <= data_col142[47];
   data_col142[49] <= data_col142[48];
   data_col142[50] <= data_col142[49];
   data_col142[51] <= data_col142[50];
   data_col142[52] <= data_col142[51];
   data_col142[53] <= data_col142[52];
   data_col142[54] <= data_col142[53];
   data_col142[55] <= data_col142[54];
   data_col142[56] <= data_col142[55];
   data_col142[57] <= data_col142[56];
   data_col142[58] <= data_col142[57];
   data_col142[59] <= data_col142[58];
   data_col142[60] <= data_col142[59];
   data_col142[61] <= data_col142[60];
   data_col142[62] <= data_col142[61];
   data_col142[63] <= data_col142[62];
   data_col142[64] <= data_col142[63];
   data_col142[65] <= data_col142[64];
   data_col142[66] <= data_col142[65];
   data_col142[67] <= data_col142[66];
   data_col142[68] <= data_col142[67];
   data_col142[69] <= data_col142[68];
   data_col142[70] <= data_col142[69];
   data_col142[71] <= data_col142[70];
   data_col142[72] <= data_col142[71];
   data_col142[73] <= data_col142[72];
   data_col142[74] <= data_col142[73];
   data_col142[75] <= data_col142[74];
   data_col142[76] <= data_col142[75];
   data_col142[77] <= data_col142[76];
   data_col142[78] <= data_col142[77];
   data_col142[79] <= data_col142[78];
   data_col142[80] <= data_col142[79];
   data_col142[81] <= data_col142[80];
   data_col142[82] <= data_col142[81];
   data_col142[83] <= data_col142[82];
   data_col142[84] <= data_col142[83];
   data_col142[85] <= data_col142[84];
   data_col142[86] <= data_col142[85];
   data_col142[87] <= data_col142[86];
   data_col142[88] <= data_col142[87];
   data_col142[89] <= data_col142[88];
   data_col142[90] <= data_col142[89];
   data_col142[91] <= data_col142[90];
   data_col142[92] <= data_col142[91];
   data_col142[93] <= data_col142[92];
   data_col142[94] <= data_col142[93];
   data_col142[95] <= data_col142[94];
   data_col142[96] <= data_col142[95];
   data_col142[97] <= data_col142[96];
   data_col142[98] <= data_col142[97];
   data_col142[99] <= data_col142[98];
   data_col142[100] <= data_col142[99];
   data_col142[101] <= data_col142[100];
   data_col142[102] <= data_col142[101];
   data_col142[103] <= data_col142[102];
   data_col142[104] <= data_col142[103];
   data_col142[105] <= data_col142[104];
   data_col142[106] <= data_col142[105];
   data_col142[107] <= data_col142[106];
   data_col142[108] <= data_col142[107];
   data_col142[109] <= data_col142[108];
   data_col142[110] <= data_col142[109];
   data_col142[111] <= data_col142[110];
   data_col142[112] <= data_col142[111];
   data_col142[113] <= data_col142[112];
   data_col142[114] <= data_col142[113];
   data_col142[115] <= data_col142[114];
   data_col142[116] <= data_col142[115];
   data_col142[117] <= data_col142[116];
   data_col142[118] <= data_col142[117];
   data_col142[119] <= data_col142[118];
   data_col142[120] <= data_col142[119];
   data_col142[121] <= data_col142[120];
   data_col142[122] <= data_col142[121];
   data_col142[123] <= data_col142[122];
   data_col142[124] <= data_col142[123];
   data_col142[125] <= data_col142[124];
   data_col142[126] <= data_col142[125];
   data_col142[127] <= data_col142[126];
   data_col142[128] <= data_col142[127];
   data_col142[129] <= data_col142[128];
   data_col142[130] <= data_col142[129];
   data_col142[131] <= data_col142[130];
   data_col142[132] <= data_col142[131];
   data_col142[133] <= data_col142[132];
   data_col142[134] <= data_col142[133];
   data_col142[135] <= data_col142[134];
   data_col142[136] <= data_col142[135];
   data_col142[137] <= data_col142[136];
   data_col142[138] <= data_col142[137];
   data_col142[139] <= data_col142[138];
   data_col142[140] <= data_col142[139];
   data_col142[141] <= data_col142[140];
   data_col142[142] <= data_col142[141];

   data_col143[1] <= data[22];
   data_col143[2] <= data_col143[1];
   data_col143[3] <= data_col143[2];
   data_col143[4] <= data_col143[3];
   data_col143[5] <= data_col143[4];
   data_col143[6] <= data_col143[5];
   data_col143[7] <= data_col143[6];
   data_col143[8] <= data_col143[7];
   data_col143[9] <= data_col143[8];
   data_col143[10] <= data_col143[9];
   data_col143[11] <= data_col143[10];
   data_col143[12] <= data_col143[11];
   data_col143[13] <= data_col143[12];
   data_col143[14] <= data_col143[13];
   data_col143[15] <= data_col143[14];
   data_col143[16] <= data_col143[15];
   data_col143[17] <= data_col143[16];
   data_col143[18] <= data_col143[17];
   data_col143[19] <= data_col143[18];
   data_col143[20] <= data_col143[19];
   data_col143[21] <= data_col143[20];
   data_col143[22] <= data_col143[21];
   data_col143[23] <= data_col143[22];
   data_col143[24] <= data_col143[23];
   data_col143[25] <= data_col143[24];
   data_col143[26] <= data_col143[25];
   data_col143[27] <= data_col143[26];
   data_col143[28] <= data_col143[27];
   data_col143[29] <= data_col143[28];
   data_col143[30] <= data_col143[29];
   data_col143[31] <= data_col143[30];
   data_col143[32] <= data_col143[31];
   data_col143[33] <= data_col143[32];
   data_col143[34] <= data_col143[33];
   data_col143[35] <= data_col143[34];
   data_col143[36] <= data_col143[35];
   data_col143[37] <= data_col143[36];
   data_col143[38] <= data_col143[37];
   data_col143[39] <= data_col143[38];
   data_col143[40] <= data_col143[39];
   data_col143[41] <= data_col143[40];
   data_col143[42] <= data_col143[41];
   data_col143[43] <= data_col143[42];
   data_col143[44] <= data_col143[43];
   data_col143[45] <= data_col143[44];
   data_col143[46] <= data_col143[45];
   data_col143[47] <= data_col143[46];
   data_col143[48] <= data_col143[47];
   data_col143[49] <= data_col143[48];
   data_col143[50] <= data_col143[49];
   data_col143[51] <= data_col143[50];
   data_col143[52] <= data_col143[51];
   data_col143[53] <= data_col143[52];
   data_col143[54] <= data_col143[53];
   data_col143[55] <= data_col143[54];
   data_col143[56] <= data_col143[55];
   data_col143[57] <= data_col143[56];
   data_col143[58] <= data_col143[57];
   data_col143[59] <= data_col143[58];
   data_col143[60] <= data_col143[59];
   data_col143[61] <= data_col143[60];
   data_col143[62] <= data_col143[61];
   data_col143[63] <= data_col143[62];
   data_col143[64] <= data_col143[63];
   data_col143[65] <= data_col143[64];
   data_col143[66] <= data_col143[65];
   data_col143[67] <= data_col143[66];
   data_col143[68] <= data_col143[67];
   data_col143[69] <= data_col143[68];
   data_col143[70] <= data_col143[69];
   data_col143[71] <= data_col143[70];
   data_col143[72] <= data_col143[71];
   data_col143[73] <= data_col143[72];
   data_col143[74] <= data_col143[73];
   data_col143[75] <= data_col143[74];
   data_col143[76] <= data_col143[75];
   data_col143[77] <= data_col143[76];
   data_col143[78] <= data_col143[77];
   data_col143[79] <= data_col143[78];
   data_col143[80] <= data_col143[79];
   data_col143[81] <= data_col143[80];
   data_col143[82] <= data_col143[81];
   data_col143[83] <= data_col143[82];
   data_col143[84] <= data_col143[83];
   data_col143[85] <= data_col143[84];
   data_col143[86] <= data_col143[85];
   data_col143[87] <= data_col143[86];
   data_col143[88] <= data_col143[87];
   data_col143[89] <= data_col143[88];
   data_col143[90] <= data_col143[89];
   data_col143[91] <= data_col143[90];
   data_col143[92] <= data_col143[91];
   data_col143[93] <= data_col143[92];
   data_col143[94] <= data_col143[93];
   data_col143[95] <= data_col143[94];
   data_col143[96] <= data_col143[95];
   data_col143[97] <= data_col143[96];
   data_col143[98] <= data_col143[97];
   data_col143[99] <= data_col143[98];
   data_col143[100] <= data_col143[99];
   data_col143[101] <= data_col143[100];
   data_col143[102] <= data_col143[101];
   data_col143[103] <= data_col143[102];
   data_col143[104] <= data_col143[103];
   data_col143[105] <= data_col143[104];
   data_col143[106] <= data_col143[105];
   data_col143[107] <= data_col143[106];
   data_col143[108] <= data_col143[107];
   data_col143[109] <= data_col143[108];
   data_col143[110] <= data_col143[109];
   data_col143[111] <= data_col143[110];
   data_col143[112] <= data_col143[111];
   data_col143[113] <= data_col143[112];
   data_col143[114] <= data_col143[113];
   data_col143[115] <= data_col143[114];
   data_col143[116] <= data_col143[115];
   data_col143[117] <= data_col143[116];
   data_col143[118] <= data_col143[117];
   data_col143[119] <= data_col143[118];
   data_col143[120] <= data_col143[119];
   data_col143[121] <= data_col143[120];
   data_col143[122] <= data_col143[121];
   data_col143[123] <= data_col143[122];
   data_col143[124] <= data_col143[123];
   data_col143[125] <= data_col143[124];
   data_col143[126] <= data_col143[125];
   data_col143[127] <= data_col143[126];
   data_col143[128] <= data_col143[127];
   data_col143[129] <= data_col143[128];
   data_col143[130] <= data_col143[129];
   data_col143[131] <= data_col143[130];
   data_col143[132] <= data_col143[131];
   data_col143[133] <= data_col143[132];
   data_col143[134] <= data_col143[133];
   data_col143[135] <= data_col143[134];
   data_col143[136] <= data_col143[135];
   data_col143[137] <= data_col143[136];
   data_col143[138] <= data_col143[137];
   data_col143[139] <= data_col143[138];
   data_col143[140] <= data_col143[139];
   data_col143[141] <= data_col143[140];
   data_col143[142] <= data_col143[141];
   data_col143[143] <= data_col143[142];

   data_col144[1] <= data[21];
   data_col144[2] <= data_col144[1];
   data_col144[3] <= data_col144[2];
   data_col144[4] <= data_col144[3];
   data_col144[5] <= data_col144[4];
   data_col144[6] <= data_col144[5];
   data_col144[7] <= data_col144[6];
   data_col144[8] <= data_col144[7];
   data_col144[9] <= data_col144[8];
   data_col144[10] <= data_col144[9];
   data_col144[11] <= data_col144[10];
   data_col144[12] <= data_col144[11];
   data_col144[13] <= data_col144[12];
   data_col144[14] <= data_col144[13];
   data_col144[15] <= data_col144[14];
   data_col144[16] <= data_col144[15];
   data_col144[17] <= data_col144[16];
   data_col144[18] <= data_col144[17];
   data_col144[19] <= data_col144[18];
   data_col144[20] <= data_col144[19];
   data_col144[21] <= data_col144[20];
   data_col144[22] <= data_col144[21];
   data_col144[23] <= data_col144[22];
   data_col144[24] <= data_col144[23];
   data_col144[25] <= data_col144[24];
   data_col144[26] <= data_col144[25];
   data_col144[27] <= data_col144[26];
   data_col144[28] <= data_col144[27];
   data_col144[29] <= data_col144[28];
   data_col144[30] <= data_col144[29];
   data_col144[31] <= data_col144[30];
   data_col144[32] <= data_col144[31];
   data_col144[33] <= data_col144[32];
   data_col144[34] <= data_col144[33];
   data_col144[35] <= data_col144[34];
   data_col144[36] <= data_col144[35];
   data_col144[37] <= data_col144[36];
   data_col144[38] <= data_col144[37];
   data_col144[39] <= data_col144[38];
   data_col144[40] <= data_col144[39];
   data_col144[41] <= data_col144[40];
   data_col144[42] <= data_col144[41];
   data_col144[43] <= data_col144[42];
   data_col144[44] <= data_col144[43];
   data_col144[45] <= data_col144[44];
   data_col144[46] <= data_col144[45];
   data_col144[47] <= data_col144[46];
   data_col144[48] <= data_col144[47];
   data_col144[49] <= data_col144[48];
   data_col144[50] <= data_col144[49];
   data_col144[51] <= data_col144[50];
   data_col144[52] <= data_col144[51];
   data_col144[53] <= data_col144[52];
   data_col144[54] <= data_col144[53];
   data_col144[55] <= data_col144[54];
   data_col144[56] <= data_col144[55];
   data_col144[57] <= data_col144[56];
   data_col144[58] <= data_col144[57];
   data_col144[59] <= data_col144[58];
   data_col144[60] <= data_col144[59];
   data_col144[61] <= data_col144[60];
   data_col144[62] <= data_col144[61];
   data_col144[63] <= data_col144[62];
   data_col144[64] <= data_col144[63];
   data_col144[65] <= data_col144[64];
   data_col144[66] <= data_col144[65];
   data_col144[67] <= data_col144[66];
   data_col144[68] <= data_col144[67];
   data_col144[69] <= data_col144[68];
   data_col144[70] <= data_col144[69];
   data_col144[71] <= data_col144[70];
   data_col144[72] <= data_col144[71];
   data_col144[73] <= data_col144[72];
   data_col144[74] <= data_col144[73];
   data_col144[75] <= data_col144[74];
   data_col144[76] <= data_col144[75];
   data_col144[77] <= data_col144[76];
   data_col144[78] <= data_col144[77];
   data_col144[79] <= data_col144[78];
   data_col144[80] <= data_col144[79];
   data_col144[81] <= data_col144[80];
   data_col144[82] <= data_col144[81];
   data_col144[83] <= data_col144[82];
   data_col144[84] <= data_col144[83];
   data_col144[85] <= data_col144[84];
   data_col144[86] <= data_col144[85];
   data_col144[87] <= data_col144[86];
   data_col144[88] <= data_col144[87];
   data_col144[89] <= data_col144[88];
   data_col144[90] <= data_col144[89];
   data_col144[91] <= data_col144[90];
   data_col144[92] <= data_col144[91];
   data_col144[93] <= data_col144[92];
   data_col144[94] <= data_col144[93];
   data_col144[95] <= data_col144[94];
   data_col144[96] <= data_col144[95];
   data_col144[97] <= data_col144[96];
   data_col144[98] <= data_col144[97];
   data_col144[99] <= data_col144[98];
   data_col144[100] <= data_col144[99];
   data_col144[101] <= data_col144[100];
   data_col144[102] <= data_col144[101];
   data_col144[103] <= data_col144[102];
   data_col144[104] <= data_col144[103];
   data_col144[105] <= data_col144[104];
   data_col144[106] <= data_col144[105];
   data_col144[107] <= data_col144[106];
   data_col144[108] <= data_col144[107];
   data_col144[109] <= data_col144[108];
   data_col144[110] <= data_col144[109];
   data_col144[111] <= data_col144[110];
   data_col144[112] <= data_col144[111];
   data_col144[113] <= data_col144[112];
   data_col144[114] <= data_col144[113];
   data_col144[115] <= data_col144[114];
   data_col144[116] <= data_col144[115];
   data_col144[117] <= data_col144[116];
   data_col144[118] <= data_col144[117];
   data_col144[119] <= data_col144[118];
   data_col144[120] <= data_col144[119];
   data_col144[121] <= data_col144[120];
   data_col144[122] <= data_col144[121];
   data_col144[123] <= data_col144[122];
   data_col144[124] <= data_col144[123];
   data_col144[125] <= data_col144[124];
   data_col144[126] <= data_col144[125];
   data_col144[127] <= data_col144[126];
   data_col144[128] <= data_col144[127];
   data_col144[129] <= data_col144[128];
   data_col144[130] <= data_col144[129];
   data_col144[131] <= data_col144[130];
   data_col144[132] <= data_col144[131];
   data_col144[133] <= data_col144[132];
   data_col144[134] <= data_col144[133];
   data_col144[135] <= data_col144[134];
   data_col144[136] <= data_col144[135];
   data_col144[137] <= data_col144[136];
   data_col144[138] <= data_col144[137];
   data_col144[139] <= data_col144[138];
   data_col144[140] <= data_col144[139];
   data_col144[141] <= data_col144[140];
   data_col144[142] <= data_col144[141];
   data_col144[143] <= data_col144[142];
   data_col144[144] <= data_col144[143];

   data_col145[1] <= data[20];
   data_col145[2] <= data_col145[1];
   data_col145[3] <= data_col145[2];
   data_col145[4] <= data_col145[3];
   data_col145[5] <= data_col145[4];
   data_col145[6] <= data_col145[5];
   data_col145[7] <= data_col145[6];
   data_col145[8] <= data_col145[7];
   data_col145[9] <= data_col145[8];
   data_col145[10] <= data_col145[9];
   data_col145[11] <= data_col145[10];
   data_col145[12] <= data_col145[11];
   data_col145[13] <= data_col145[12];
   data_col145[14] <= data_col145[13];
   data_col145[15] <= data_col145[14];
   data_col145[16] <= data_col145[15];
   data_col145[17] <= data_col145[16];
   data_col145[18] <= data_col145[17];
   data_col145[19] <= data_col145[18];
   data_col145[20] <= data_col145[19];
   data_col145[21] <= data_col145[20];
   data_col145[22] <= data_col145[21];
   data_col145[23] <= data_col145[22];
   data_col145[24] <= data_col145[23];
   data_col145[25] <= data_col145[24];
   data_col145[26] <= data_col145[25];
   data_col145[27] <= data_col145[26];
   data_col145[28] <= data_col145[27];
   data_col145[29] <= data_col145[28];
   data_col145[30] <= data_col145[29];
   data_col145[31] <= data_col145[30];
   data_col145[32] <= data_col145[31];
   data_col145[33] <= data_col145[32];
   data_col145[34] <= data_col145[33];
   data_col145[35] <= data_col145[34];
   data_col145[36] <= data_col145[35];
   data_col145[37] <= data_col145[36];
   data_col145[38] <= data_col145[37];
   data_col145[39] <= data_col145[38];
   data_col145[40] <= data_col145[39];
   data_col145[41] <= data_col145[40];
   data_col145[42] <= data_col145[41];
   data_col145[43] <= data_col145[42];
   data_col145[44] <= data_col145[43];
   data_col145[45] <= data_col145[44];
   data_col145[46] <= data_col145[45];
   data_col145[47] <= data_col145[46];
   data_col145[48] <= data_col145[47];
   data_col145[49] <= data_col145[48];
   data_col145[50] <= data_col145[49];
   data_col145[51] <= data_col145[50];
   data_col145[52] <= data_col145[51];
   data_col145[53] <= data_col145[52];
   data_col145[54] <= data_col145[53];
   data_col145[55] <= data_col145[54];
   data_col145[56] <= data_col145[55];
   data_col145[57] <= data_col145[56];
   data_col145[58] <= data_col145[57];
   data_col145[59] <= data_col145[58];
   data_col145[60] <= data_col145[59];
   data_col145[61] <= data_col145[60];
   data_col145[62] <= data_col145[61];
   data_col145[63] <= data_col145[62];
   data_col145[64] <= data_col145[63];
   data_col145[65] <= data_col145[64];
   data_col145[66] <= data_col145[65];
   data_col145[67] <= data_col145[66];
   data_col145[68] <= data_col145[67];
   data_col145[69] <= data_col145[68];
   data_col145[70] <= data_col145[69];
   data_col145[71] <= data_col145[70];
   data_col145[72] <= data_col145[71];
   data_col145[73] <= data_col145[72];
   data_col145[74] <= data_col145[73];
   data_col145[75] <= data_col145[74];
   data_col145[76] <= data_col145[75];
   data_col145[77] <= data_col145[76];
   data_col145[78] <= data_col145[77];
   data_col145[79] <= data_col145[78];
   data_col145[80] <= data_col145[79];
   data_col145[81] <= data_col145[80];
   data_col145[82] <= data_col145[81];
   data_col145[83] <= data_col145[82];
   data_col145[84] <= data_col145[83];
   data_col145[85] <= data_col145[84];
   data_col145[86] <= data_col145[85];
   data_col145[87] <= data_col145[86];
   data_col145[88] <= data_col145[87];
   data_col145[89] <= data_col145[88];
   data_col145[90] <= data_col145[89];
   data_col145[91] <= data_col145[90];
   data_col145[92] <= data_col145[91];
   data_col145[93] <= data_col145[92];
   data_col145[94] <= data_col145[93];
   data_col145[95] <= data_col145[94];
   data_col145[96] <= data_col145[95];
   data_col145[97] <= data_col145[96];
   data_col145[98] <= data_col145[97];
   data_col145[99] <= data_col145[98];
   data_col145[100] <= data_col145[99];
   data_col145[101] <= data_col145[100];
   data_col145[102] <= data_col145[101];
   data_col145[103] <= data_col145[102];
   data_col145[104] <= data_col145[103];
   data_col145[105] <= data_col145[104];
   data_col145[106] <= data_col145[105];
   data_col145[107] <= data_col145[106];
   data_col145[108] <= data_col145[107];
   data_col145[109] <= data_col145[108];
   data_col145[110] <= data_col145[109];
   data_col145[111] <= data_col145[110];
   data_col145[112] <= data_col145[111];
   data_col145[113] <= data_col145[112];
   data_col145[114] <= data_col145[113];
   data_col145[115] <= data_col145[114];
   data_col145[116] <= data_col145[115];
   data_col145[117] <= data_col145[116];
   data_col145[118] <= data_col145[117];
   data_col145[119] <= data_col145[118];
   data_col145[120] <= data_col145[119];
   data_col145[121] <= data_col145[120];
   data_col145[122] <= data_col145[121];
   data_col145[123] <= data_col145[122];
   data_col145[124] <= data_col145[123];
   data_col145[125] <= data_col145[124];
   data_col145[126] <= data_col145[125];
   data_col145[127] <= data_col145[126];
   data_col145[128] <= data_col145[127];
   data_col145[129] <= data_col145[128];
   data_col145[130] <= data_col145[129];
   data_col145[131] <= data_col145[130];
   data_col145[132] <= data_col145[131];
   data_col145[133] <= data_col145[132];
   data_col145[134] <= data_col145[133];
   data_col145[135] <= data_col145[134];
   data_col145[136] <= data_col145[135];
   data_col145[137] <= data_col145[136];
   data_col145[138] <= data_col145[137];
   data_col145[139] <= data_col145[138];
   data_col145[140] <= data_col145[139];
   data_col145[141] <= data_col145[140];
   data_col145[142] <= data_col145[141];
   data_col145[143] <= data_col145[142];
   data_col145[144] <= data_col145[143];
   data_col145[145] <= data_col145[144];

   data_col146[1] <= data[19];
   data_col146[2] <= data_col146[1];
   data_col146[3] <= data_col146[2];
   data_col146[4] <= data_col146[3];
   data_col146[5] <= data_col146[4];
   data_col146[6] <= data_col146[5];
   data_col146[7] <= data_col146[6];
   data_col146[8] <= data_col146[7];
   data_col146[9] <= data_col146[8];
   data_col146[10] <= data_col146[9];
   data_col146[11] <= data_col146[10];
   data_col146[12] <= data_col146[11];
   data_col146[13] <= data_col146[12];
   data_col146[14] <= data_col146[13];
   data_col146[15] <= data_col146[14];
   data_col146[16] <= data_col146[15];
   data_col146[17] <= data_col146[16];
   data_col146[18] <= data_col146[17];
   data_col146[19] <= data_col146[18];
   data_col146[20] <= data_col146[19];
   data_col146[21] <= data_col146[20];
   data_col146[22] <= data_col146[21];
   data_col146[23] <= data_col146[22];
   data_col146[24] <= data_col146[23];
   data_col146[25] <= data_col146[24];
   data_col146[26] <= data_col146[25];
   data_col146[27] <= data_col146[26];
   data_col146[28] <= data_col146[27];
   data_col146[29] <= data_col146[28];
   data_col146[30] <= data_col146[29];
   data_col146[31] <= data_col146[30];
   data_col146[32] <= data_col146[31];
   data_col146[33] <= data_col146[32];
   data_col146[34] <= data_col146[33];
   data_col146[35] <= data_col146[34];
   data_col146[36] <= data_col146[35];
   data_col146[37] <= data_col146[36];
   data_col146[38] <= data_col146[37];
   data_col146[39] <= data_col146[38];
   data_col146[40] <= data_col146[39];
   data_col146[41] <= data_col146[40];
   data_col146[42] <= data_col146[41];
   data_col146[43] <= data_col146[42];
   data_col146[44] <= data_col146[43];
   data_col146[45] <= data_col146[44];
   data_col146[46] <= data_col146[45];
   data_col146[47] <= data_col146[46];
   data_col146[48] <= data_col146[47];
   data_col146[49] <= data_col146[48];
   data_col146[50] <= data_col146[49];
   data_col146[51] <= data_col146[50];
   data_col146[52] <= data_col146[51];
   data_col146[53] <= data_col146[52];
   data_col146[54] <= data_col146[53];
   data_col146[55] <= data_col146[54];
   data_col146[56] <= data_col146[55];
   data_col146[57] <= data_col146[56];
   data_col146[58] <= data_col146[57];
   data_col146[59] <= data_col146[58];
   data_col146[60] <= data_col146[59];
   data_col146[61] <= data_col146[60];
   data_col146[62] <= data_col146[61];
   data_col146[63] <= data_col146[62];
   data_col146[64] <= data_col146[63];
   data_col146[65] <= data_col146[64];
   data_col146[66] <= data_col146[65];
   data_col146[67] <= data_col146[66];
   data_col146[68] <= data_col146[67];
   data_col146[69] <= data_col146[68];
   data_col146[70] <= data_col146[69];
   data_col146[71] <= data_col146[70];
   data_col146[72] <= data_col146[71];
   data_col146[73] <= data_col146[72];
   data_col146[74] <= data_col146[73];
   data_col146[75] <= data_col146[74];
   data_col146[76] <= data_col146[75];
   data_col146[77] <= data_col146[76];
   data_col146[78] <= data_col146[77];
   data_col146[79] <= data_col146[78];
   data_col146[80] <= data_col146[79];
   data_col146[81] <= data_col146[80];
   data_col146[82] <= data_col146[81];
   data_col146[83] <= data_col146[82];
   data_col146[84] <= data_col146[83];
   data_col146[85] <= data_col146[84];
   data_col146[86] <= data_col146[85];
   data_col146[87] <= data_col146[86];
   data_col146[88] <= data_col146[87];
   data_col146[89] <= data_col146[88];
   data_col146[90] <= data_col146[89];
   data_col146[91] <= data_col146[90];
   data_col146[92] <= data_col146[91];
   data_col146[93] <= data_col146[92];
   data_col146[94] <= data_col146[93];
   data_col146[95] <= data_col146[94];
   data_col146[96] <= data_col146[95];
   data_col146[97] <= data_col146[96];
   data_col146[98] <= data_col146[97];
   data_col146[99] <= data_col146[98];
   data_col146[100] <= data_col146[99];
   data_col146[101] <= data_col146[100];
   data_col146[102] <= data_col146[101];
   data_col146[103] <= data_col146[102];
   data_col146[104] <= data_col146[103];
   data_col146[105] <= data_col146[104];
   data_col146[106] <= data_col146[105];
   data_col146[107] <= data_col146[106];
   data_col146[108] <= data_col146[107];
   data_col146[109] <= data_col146[108];
   data_col146[110] <= data_col146[109];
   data_col146[111] <= data_col146[110];
   data_col146[112] <= data_col146[111];
   data_col146[113] <= data_col146[112];
   data_col146[114] <= data_col146[113];
   data_col146[115] <= data_col146[114];
   data_col146[116] <= data_col146[115];
   data_col146[117] <= data_col146[116];
   data_col146[118] <= data_col146[117];
   data_col146[119] <= data_col146[118];
   data_col146[120] <= data_col146[119];
   data_col146[121] <= data_col146[120];
   data_col146[122] <= data_col146[121];
   data_col146[123] <= data_col146[122];
   data_col146[124] <= data_col146[123];
   data_col146[125] <= data_col146[124];
   data_col146[126] <= data_col146[125];
   data_col146[127] <= data_col146[126];
   data_col146[128] <= data_col146[127];
   data_col146[129] <= data_col146[128];
   data_col146[130] <= data_col146[129];
   data_col146[131] <= data_col146[130];
   data_col146[132] <= data_col146[131];
   data_col146[133] <= data_col146[132];
   data_col146[134] <= data_col146[133];
   data_col146[135] <= data_col146[134];
   data_col146[136] <= data_col146[135];
   data_col146[137] <= data_col146[136];
   data_col146[138] <= data_col146[137];
   data_col146[139] <= data_col146[138];
   data_col146[140] <= data_col146[139];
   data_col146[141] <= data_col146[140];
   data_col146[142] <= data_col146[141];
   data_col146[143] <= data_col146[142];
   data_col146[144] <= data_col146[143];
   data_col146[145] <= data_col146[144];
   data_col146[146] <= data_col146[145];

   data_col147[1] <= data[18];
   data_col147[2] <= data_col147[1];
   data_col147[3] <= data_col147[2];
   data_col147[4] <= data_col147[3];
   data_col147[5] <= data_col147[4];
   data_col147[6] <= data_col147[5];
   data_col147[7] <= data_col147[6];
   data_col147[8] <= data_col147[7];
   data_col147[9] <= data_col147[8];
   data_col147[10] <= data_col147[9];
   data_col147[11] <= data_col147[10];
   data_col147[12] <= data_col147[11];
   data_col147[13] <= data_col147[12];
   data_col147[14] <= data_col147[13];
   data_col147[15] <= data_col147[14];
   data_col147[16] <= data_col147[15];
   data_col147[17] <= data_col147[16];
   data_col147[18] <= data_col147[17];
   data_col147[19] <= data_col147[18];
   data_col147[20] <= data_col147[19];
   data_col147[21] <= data_col147[20];
   data_col147[22] <= data_col147[21];
   data_col147[23] <= data_col147[22];
   data_col147[24] <= data_col147[23];
   data_col147[25] <= data_col147[24];
   data_col147[26] <= data_col147[25];
   data_col147[27] <= data_col147[26];
   data_col147[28] <= data_col147[27];
   data_col147[29] <= data_col147[28];
   data_col147[30] <= data_col147[29];
   data_col147[31] <= data_col147[30];
   data_col147[32] <= data_col147[31];
   data_col147[33] <= data_col147[32];
   data_col147[34] <= data_col147[33];
   data_col147[35] <= data_col147[34];
   data_col147[36] <= data_col147[35];
   data_col147[37] <= data_col147[36];
   data_col147[38] <= data_col147[37];
   data_col147[39] <= data_col147[38];
   data_col147[40] <= data_col147[39];
   data_col147[41] <= data_col147[40];
   data_col147[42] <= data_col147[41];
   data_col147[43] <= data_col147[42];
   data_col147[44] <= data_col147[43];
   data_col147[45] <= data_col147[44];
   data_col147[46] <= data_col147[45];
   data_col147[47] <= data_col147[46];
   data_col147[48] <= data_col147[47];
   data_col147[49] <= data_col147[48];
   data_col147[50] <= data_col147[49];
   data_col147[51] <= data_col147[50];
   data_col147[52] <= data_col147[51];
   data_col147[53] <= data_col147[52];
   data_col147[54] <= data_col147[53];
   data_col147[55] <= data_col147[54];
   data_col147[56] <= data_col147[55];
   data_col147[57] <= data_col147[56];
   data_col147[58] <= data_col147[57];
   data_col147[59] <= data_col147[58];
   data_col147[60] <= data_col147[59];
   data_col147[61] <= data_col147[60];
   data_col147[62] <= data_col147[61];
   data_col147[63] <= data_col147[62];
   data_col147[64] <= data_col147[63];
   data_col147[65] <= data_col147[64];
   data_col147[66] <= data_col147[65];
   data_col147[67] <= data_col147[66];
   data_col147[68] <= data_col147[67];
   data_col147[69] <= data_col147[68];
   data_col147[70] <= data_col147[69];
   data_col147[71] <= data_col147[70];
   data_col147[72] <= data_col147[71];
   data_col147[73] <= data_col147[72];
   data_col147[74] <= data_col147[73];
   data_col147[75] <= data_col147[74];
   data_col147[76] <= data_col147[75];
   data_col147[77] <= data_col147[76];
   data_col147[78] <= data_col147[77];
   data_col147[79] <= data_col147[78];
   data_col147[80] <= data_col147[79];
   data_col147[81] <= data_col147[80];
   data_col147[82] <= data_col147[81];
   data_col147[83] <= data_col147[82];
   data_col147[84] <= data_col147[83];
   data_col147[85] <= data_col147[84];
   data_col147[86] <= data_col147[85];
   data_col147[87] <= data_col147[86];
   data_col147[88] <= data_col147[87];
   data_col147[89] <= data_col147[88];
   data_col147[90] <= data_col147[89];
   data_col147[91] <= data_col147[90];
   data_col147[92] <= data_col147[91];
   data_col147[93] <= data_col147[92];
   data_col147[94] <= data_col147[93];
   data_col147[95] <= data_col147[94];
   data_col147[96] <= data_col147[95];
   data_col147[97] <= data_col147[96];
   data_col147[98] <= data_col147[97];
   data_col147[99] <= data_col147[98];
   data_col147[100] <= data_col147[99];
   data_col147[101] <= data_col147[100];
   data_col147[102] <= data_col147[101];
   data_col147[103] <= data_col147[102];
   data_col147[104] <= data_col147[103];
   data_col147[105] <= data_col147[104];
   data_col147[106] <= data_col147[105];
   data_col147[107] <= data_col147[106];
   data_col147[108] <= data_col147[107];
   data_col147[109] <= data_col147[108];
   data_col147[110] <= data_col147[109];
   data_col147[111] <= data_col147[110];
   data_col147[112] <= data_col147[111];
   data_col147[113] <= data_col147[112];
   data_col147[114] <= data_col147[113];
   data_col147[115] <= data_col147[114];
   data_col147[116] <= data_col147[115];
   data_col147[117] <= data_col147[116];
   data_col147[118] <= data_col147[117];
   data_col147[119] <= data_col147[118];
   data_col147[120] <= data_col147[119];
   data_col147[121] <= data_col147[120];
   data_col147[122] <= data_col147[121];
   data_col147[123] <= data_col147[122];
   data_col147[124] <= data_col147[123];
   data_col147[125] <= data_col147[124];
   data_col147[126] <= data_col147[125];
   data_col147[127] <= data_col147[126];
   data_col147[128] <= data_col147[127];
   data_col147[129] <= data_col147[128];
   data_col147[130] <= data_col147[129];
   data_col147[131] <= data_col147[130];
   data_col147[132] <= data_col147[131];
   data_col147[133] <= data_col147[132];
   data_col147[134] <= data_col147[133];
   data_col147[135] <= data_col147[134];
   data_col147[136] <= data_col147[135];
   data_col147[137] <= data_col147[136];
   data_col147[138] <= data_col147[137];
   data_col147[139] <= data_col147[138];
   data_col147[140] <= data_col147[139];
   data_col147[141] <= data_col147[140];
   data_col147[142] <= data_col147[141];
   data_col147[143] <= data_col147[142];
   data_col147[144] <= data_col147[143];
   data_col147[145] <= data_col147[144];
   data_col147[146] <= data_col147[145];
   data_col147[147] <= data_col147[146];

   data_col148[1] <= data[17];
   data_col148[2] <= data_col148[1];
   data_col148[3] <= data_col148[2];
   data_col148[4] <= data_col148[3];
   data_col148[5] <= data_col148[4];
   data_col148[6] <= data_col148[5];
   data_col148[7] <= data_col148[6];
   data_col148[8] <= data_col148[7];
   data_col148[9] <= data_col148[8];
   data_col148[10] <= data_col148[9];
   data_col148[11] <= data_col148[10];
   data_col148[12] <= data_col148[11];
   data_col148[13] <= data_col148[12];
   data_col148[14] <= data_col148[13];
   data_col148[15] <= data_col148[14];
   data_col148[16] <= data_col148[15];
   data_col148[17] <= data_col148[16];
   data_col148[18] <= data_col148[17];
   data_col148[19] <= data_col148[18];
   data_col148[20] <= data_col148[19];
   data_col148[21] <= data_col148[20];
   data_col148[22] <= data_col148[21];
   data_col148[23] <= data_col148[22];
   data_col148[24] <= data_col148[23];
   data_col148[25] <= data_col148[24];
   data_col148[26] <= data_col148[25];
   data_col148[27] <= data_col148[26];
   data_col148[28] <= data_col148[27];
   data_col148[29] <= data_col148[28];
   data_col148[30] <= data_col148[29];
   data_col148[31] <= data_col148[30];
   data_col148[32] <= data_col148[31];
   data_col148[33] <= data_col148[32];
   data_col148[34] <= data_col148[33];
   data_col148[35] <= data_col148[34];
   data_col148[36] <= data_col148[35];
   data_col148[37] <= data_col148[36];
   data_col148[38] <= data_col148[37];
   data_col148[39] <= data_col148[38];
   data_col148[40] <= data_col148[39];
   data_col148[41] <= data_col148[40];
   data_col148[42] <= data_col148[41];
   data_col148[43] <= data_col148[42];
   data_col148[44] <= data_col148[43];
   data_col148[45] <= data_col148[44];
   data_col148[46] <= data_col148[45];
   data_col148[47] <= data_col148[46];
   data_col148[48] <= data_col148[47];
   data_col148[49] <= data_col148[48];
   data_col148[50] <= data_col148[49];
   data_col148[51] <= data_col148[50];
   data_col148[52] <= data_col148[51];
   data_col148[53] <= data_col148[52];
   data_col148[54] <= data_col148[53];
   data_col148[55] <= data_col148[54];
   data_col148[56] <= data_col148[55];
   data_col148[57] <= data_col148[56];
   data_col148[58] <= data_col148[57];
   data_col148[59] <= data_col148[58];
   data_col148[60] <= data_col148[59];
   data_col148[61] <= data_col148[60];
   data_col148[62] <= data_col148[61];
   data_col148[63] <= data_col148[62];
   data_col148[64] <= data_col148[63];
   data_col148[65] <= data_col148[64];
   data_col148[66] <= data_col148[65];
   data_col148[67] <= data_col148[66];
   data_col148[68] <= data_col148[67];
   data_col148[69] <= data_col148[68];
   data_col148[70] <= data_col148[69];
   data_col148[71] <= data_col148[70];
   data_col148[72] <= data_col148[71];
   data_col148[73] <= data_col148[72];
   data_col148[74] <= data_col148[73];
   data_col148[75] <= data_col148[74];
   data_col148[76] <= data_col148[75];
   data_col148[77] <= data_col148[76];
   data_col148[78] <= data_col148[77];
   data_col148[79] <= data_col148[78];
   data_col148[80] <= data_col148[79];
   data_col148[81] <= data_col148[80];
   data_col148[82] <= data_col148[81];
   data_col148[83] <= data_col148[82];
   data_col148[84] <= data_col148[83];
   data_col148[85] <= data_col148[84];
   data_col148[86] <= data_col148[85];
   data_col148[87] <= data_col148[86];
   data_col148[88] <= data_col148[87];
   data_col148[89] <= data_col148[88];
   data_col148[90] <= data_col148[89];
   data_col148[91] <= data_col148[90];
   data_col148[92] <= data_col148[91];
   data_col148[93] <= data_col148[92];
   data_col148[94] <= data_col148[93];
   data_col148[95] <= data_col148[94];
   data_col148[96] <= data_col148[95];
   data_col148[97] <= data_col148[96];
   data_col148[98] <= data_col148[97];
   data_col148[99] <= data_col148[98];
   data_col148[100] <= data_col148[99];
   data_col148[101] <= data_col148[100];
   data_col148[102] <= data_col148[101];
   data_col148[103] <= data_col148[102];
   data_col148[104] <= data_col148[103];
   data_col148[105] <= data_col148[104];
   data_col148[106] <= data_col148[105];
   data_col148[107] <= data_col148[106];
   data_col148[108] <= data_col148[107];
   data_col148[109] <= data_col148[108];
   data_col148[110] <= data_col148[109];
   data_col148[111] <= data_col148[110];
   data_col148[112] <= data_col148[111];
   data_col148[113] <= data_col148[112];
   data_col148[114] <= data_col148[113];
   data_col148[115] <= data_col148[114];
   data_col148[116] <= data_col148[115];
   data_col148[117] <= data_col148[116];
   data_col148[118] <= data_col148[117];
   data_col148[119] <= data_col148[118];
   data_col148[120] <= data_col148[119];
   data_col148[121] <= data_col148[120];
   data_col148[122] <= data_col148[121];
   data_col148[123] <= data_col148[122];
   data_col148[124] <= data_col148[123];
   data_col148[125] <= data_col148[124];
   data_col148[126] <= data_col148[125];
   data_col148[127] <= data_col148[126];
   data_col148[128] <= data_col148[127];
   data_col148[129] <= data_col148[128];
   data_col148[130] <= data_col148[129];
   data_col148[131] <= data_col148[130];
   data_col148[132] <= data_col148[131];
   data_col148[133] <= data_col148[132];
   data_col148[134] <= data_col148[133];
   data_col148[135] <= data_col148[134];
   data_col148[136] <= data_col148[135];
   data_col148[137] <= data_col148[136];
   data_col148[138] <= data_col148[137];
   data_col148[139] <= data_col148[138];
   data_col148[140] <= data_col148[139];
   data_col148[141] <= data_col148[140];
   data_col148[142] <= data_col148[141];
   data_col148[143] <= data_col148[142];
   data_col148[144] <= data_col148[143];
   data_col148[145] <= data_col148[144];
   data_col148[146] <= data_col148[145];
   data_col148[147] <= data_col148[146];
   data_col148[148] <= data_col148[147];

   data_col149[1] <= data[16];
   data_col149[2] <= data_col149[1];
   data_col149[3] <= data_col149[2];
   data_col149[4] <= data_col149[3];
   data_col149[5] <= data_col149[4];
   data_col149[6] <= data_col149[5];
   data_col149[7] <= data_col149[6];
   data_col149[8] <= data_col149[7];
   data_col149[9] <= data_col149[8];
   data_col149[10] <= data_col149[9];
   data_col149[11] <= data_col149[10];
   data_col149[12] <= data_col149[11];
   data_col149[13] <= data_col149[12];
   data_col149[14] <= data_col149[13];
   data_col149[15] <= data_col149[14];
   data_col149[16] <= data_col149[15];
   data_col149[17] <= data_col149[16];
   data_col149[18] <= data_col149[17];
   data_col149[19] <= data_col149[18];
   data_col149[20] <= data_col149[19];
   data_col149[21] <= data_col149[20];
   data_col149[22] <= data_col149[21];
   data_col149[23] <= data_col149[22];
   data_col149[24] <= data_col149[23];
   data_col149[25] <= data_col149[24];
   data_col149[26] <= data_col149[25];
   data_col149[27] <= data_col149[26];
   data_col149[28] <= data_col149[27];
   data_col149[29] <= data_col149[28];
   data_col149[30] <= data_col149[29];
   data_col149[31] <= data_col149[30];
   data_col149[32] <= data_col149[31];
   data_col149[33] <= data_col149[32];
   data_col149[34] <= data_col149[33];
   data_col149[35] <= data_col149[34];
   data_col149[36] <= data_col149[35];
   data_col149[37] <= data_col149[36];
   data_col149[38] <= data_col149[37];
   data_col149[39] <= data_col149[38];
   data_col149[40] <= data_col149[39];
   data_col149[41] <= data_col149[40];
   data_col149[42] <= data_col149[41];
   data_col149[43] <= data_col149[42];
   data_col149[44] <= data_col149[43];
   data_col149[45] <= data_col149[44];
   data_col149[46] <= data_col149[45];
   data_col149[47] <= data_col149[46];
   data_col149[48] <= data_col149[47];
   data_col149[49] <= data_col149[48];
   data_col149[50] <= data_col149[49];
   data_col149[51] <= data_col149[50];
   data_col149[52] <= data_col149[51];
   data_col149[53] <= data_col149[52];
   data_col149[54] <= data_col149[53];
   data_col149[55] <= data_col149[54];
   data_col149[56] <= data_col149[55];
   data_col149[57] <= data_col149[56];
   data_col149[58] <= data_col149[57];
   data_col149[59] <= data_col149[58];
   data_col149[60] <= data_col149[59];
   data_col149[61] <= data_col149[60];
   data_col149[62] <= data_col149[61];
   data_col149[63] <= data_col149[62];
   data_col149[64] <= data_col149[63];
   data_col149[65] <= data_col149[64];
   data_col149[66] <= data_col149[65];
   data_col149[67] <= data_col149[66];
   data_col149[68] <= data_col149[67];
   data_col149[69] <= data_col149[68];
   data_col149[70] <= data_col149[69];
   data_col149[71] <= data_col149[70];
   data_col149[72] <= data_col149[71];
   data_col149[73] <= data_col149[72];
   data_col149[74] <= data_col149[73];
   data_col149[75] <= data_col149[74];
   data_col149[76] <= data_col149[75];
   data_col149[77] <= data_col149[76];
   data_col149[78] <= data_col149[77];
   data_col149[79] <= data_col149[78];
   data_col149[80] <= data_col149[79];
   data_col149[81] <= data_col149[80];
   data_col149[82] <= data_col149[81];
   data_col149[83] <= data_col149[82];
   data_col149[84] <= data_col149[83];
   data_col149[85] <= data_col149[84];
   data_col149[86] <= data_col149[85];
   data_col149[87] <= data_col149[86];
   data_col149[88] <= data_col149[87];
   data_col149[89] <= data_col149[88];
   data_col149[90] <= data_col149[89];
   data_col149[91] <= data_col149[90];
   data_col149[92] <= data_col149[91];
   data_col149[93] <= data_col149[92];
   data_col149[94] <= data_col149[93];
   data_col149[95] <= data_col149[94];
   data_col149[96] <= data_col149[95];
   data_col149[97] <= data_col149[96];
   data_col149[98] <= data_col149[97];
   data_col149[99] <= data_col149[98];
   data_col149[100] <= data_col149[99];
   data_col149[101] <= data_col149[100];
   data_col149[102] <= data_col149[101];
   data_col149[103] <= data_col149[102];
   data_col149[104] <= data_col149[103];
   data_col149[105] <= data_col149[104];
   data_col149[106] <= data_col149[105];
   data_col149[107] <= data_col149[106];
   data_col149[108] <= data_col149[107];
   data_col149[109] <= data_col149[108];
   data_col149[110] <= data_col149[109];
   data_col149[111] <= data_col149[110];
   data_col149[112] <= data_col149[111];
   data_col149[113] <= data_col149[112];
   data_col149[114] <= data_col149[113];
   data_col149[115] <= data_col149[114];
   data_col149[116] <= data_col149[115];
   data_col149[117] <= data_col149[116];
   data_col149[118] <= data_col149[117];
   data_col149[119] <= data_col149[118];
   data_col149[120] <= data_col149[119];
   data_col149[121] <= data_col149[120];
   data_col149[122] <= data_col149[121];
   data_col149[123] <= data_col149[122];
   data_col149[124] <= data_col149[123];
   data_col149[125] <= data_col149[124];
   data_col149[126] <= data_col149[125];
   data_col149[127] <= data_col149[126];
   data_col149[128] <= data_col149[127];
   data_col149[129] <= data_col149[128];
   data_col149[130] <= data_col149[129];
   data_col149[131] <= data_col149[130];
   data_col149[132] <= data_col149[131];
   data_col149[133] <= data_col149[132];
   data_col149[134] <= data_col149[133];
   data_col149[135] <= data_col149[134];
   data_col149[136] <= data_col149[135];
   data_col149[137] <= data_col149[136];
   data_col149[138] <= data_col149[137];
   data_col149[139] <= data_col149[138];
   data_col149[140] <= data_col149[139];
   data_col149[141] <= data_col149[140];
   data_col149[142] <= data_col149[141];
   data_col149[143] <= data_col149[142];
   data_col149[144] <= data_col149[143];
   data_col149[145] <= data_col149[144];
   data_col149[146] <= data_col149[145];
   data_col149[147] <= data_col149[146];
   data_col149[148] <= data_col149[147];
   data_col149[149] <= data_col149[148];

   data_col150[1] <= data[15];
   data_col150[2] <= data_col150[1];
   data_col150[3] <= data_col150[2];
   data_col150[4] <= data_col150[3];
   data_col150[5] <= data_col150[4];
   data_col150[6] <= data_col150[5];
   data_col150[7] <= data_col150[6];
   data_col150[8] <= data_col150[7];
   data_col150[9] <= data_col150[8];
   data_col150[10] <= data_col150[9];
   data_col150[11] <= data_col150[10];
   data_col150[12] <= data_col150[11];
   data_col150[13] <= data_col150[12];
   data_col150[14] <= data_col150[13];
   data_col150[15] <= data_col150[14];
   data_col150[16] <= data_col150[15];
   data_col150[17] <= data_col150[16];
   data_col150[18] <= data_col150[17];
   data_col150[19] <= data_col150[18];
   data_col150[20] <= data_col150[19];
   data_col150[21] <= data_col150[20];
   data_col150[22] <= data_col150[21];
   data_col150[23] <= data_col150[22];
   data_col150[24] <= data_col150[23];
   data_col150[25] <= data_col150[24];
   data_col150[26] <= data_col150[25];
   data_col150[27] <= data_col150[26];
   data_col150[28] <= data_col150[27];
   data_col150[29] <= data_col150[28];
   data_col150[30] <= data_col150[29];
   data_col150[31] <= data_col150[30];
   data_col150[32] <= data_col150[31];
   data_col150[33] <= data_col150[32];
   data_col150[34] <= data_col150[33];
   data_col150[35] <= data_col150[34];
   data_col150[36] <= data_col150[35];
   data_col150[37] <= data_col150[36];
   data_col150[38] <= data_col150[37];
   data_col150[39] <= data_col150[38];
   data_col150[40] <= data_col150[39];
   data_col150[41] <= data_col150[40];
   data_col150[42] <= data_col150[41];
   data_col150[43] <= data_col150[42];
   data_col150[44] <= data_col150[43];
   data_col150[45] <= data_col150[44];
   data_col150[46] <= data_col150[45];
   data_col150[47] <= data_col150[46];
   data_col150[48] <= data_col150[47];
   data_col150[49] <= data_col150[48];
   data_col150[50] <= data_col150[49];
   data_col150[51] <= data_col150[50];
   data_col150[52] <= data_col150[51];
   data_col150[53] <= data_col150[52];
   data_col150[54] <= data_col150[53];
   data_col150[55] <= data_col150[54];
   data_col150[56] <= data_col150[55];
   data_col150[57] <= data_col150[56];
   data_col150[58] <= data_col150[57];
   data_col150[59] <= data_col150[58];
   data_col150[60] <= data_col150[59];
   data_col150[61] <= data_col150[60];
   data_col150[62] <= data_col150[61];
   data_col150[63] <= data_col150[62];
   data_col150[64] <= data_col150[63];
   data_col150[65] <= data_col150[64];
   data_col150[66] <= data_col150[65];
   data_col150[67] <= data_col150[66];
   data_col150[68] <= data_col150[67];
   data_col150[69] <= data_col150[68];
   data_col150[70] <= data_col150[69];
   data_col150[71] <= data_col150[70];
   data_col150[72] <= data_col150[71];
   data_col150[73] <= data_col150[72];
   data_col150[74] <= data_col150[73];
   data_col150[75] <= data_col150[74];
   data_col150[76] <= data_col150[75];
   data_col150[77] <= data_col150[76];
   data_col150[78] <= data_col150[77];
   data_col150[79] <= data_col150[78];
   data_col150[80] <= data_col150[79];
   data_col150[81] <= data_col150[80];
   data_col150[82] <= data_col150[81];
   data_col150[83] <= data_col150[82];
   data_col150[84] <= data_col150[83];
   data_col150[85] <= data_col150[84];
   data_col150[86] <= data_col150[85];
   data_col150[87] <= data_col150[86];
   data_col150[88] <= data_col150[87];
   data_col150[89] <= data_col150[88];
   data_col150[90] <= data_col150[89];
   data_col150[91] <= data_col150[90];
   data_col150[92] <= data_col150[91];
   data_col150[93] <= data_col150[92];
   data_col150[94] <= data_col150[93];
   data_col150[95] <= data_col150[94];
   data_col150[96] <= data_col150[95];
   data_col150[97] <= data_col150[96];
   data_col150[98] <= data_col150[97];
   data_col150[99] <= data_col150[98];
   data_col150[100] <= data_col150[99];
   data_col150[101] <= data_col150[100];
   data_col150[102] <= data_col150[101];
   data_col150[103] <= data_col150[102];
   data_col150[104] <= data_col150[103];
   data_col150[105] <= data_col150[104];
   data_col150[106] <= data_col150[105];
   data_col150[107] <= data_col150[106];
   data_col150[108] <= data_col150[107];
   data_col150[109] <= data_col150[108];
   data_col150[110] <= data_col150[109];
   data_col150[111] <= data_col150[110];
   data_col150[112] <= data_col150[111];
   data_col150[113] <= data_col150[112];
   data_col150[114] <= data_col150[113];
   data_col150[115] <= data_col150[114];
   data_col150[116] <= data_col150[115];
   data_col150[117] <= data_col150[116];
   data_col150[118] <= data_col150[117];
   data_col150[119] <= data_col150[118];
   data_col150[120] <= data_col150[119];
   data_col150[121] <= data_col150[120];
   data_col150[122] <= data_col150[121];
   data_col150[123] <= data_col150[122];
   data_col150[124] <= data_col150[123];
   data_col150[125] <= data_col150[124];
   data_col150[126] <= data_col150[125];
   data_col150[127] <= data_col150[126];
   data_col150[128] <= data_col150[127];
   data_col150[129] <= data_col150[128];
   data_col150[130] <= data_col150[129];
   data_col150[131] <= data_col150[130];
   data_col150[132] <= data_col150[131];
   data_col150[133] <= data_col150[132];
   data_col150[134] <= data_col150[133];
   data_col150[135] <= data_col150[134];
   data_col150[136] <= data_col150[135];
   data_col150[137] <= data_col150[136];
   data_col150[138] <= data_col150[137];
   data_col150[139] <= data_col150[138];
   data_col150[140] <= data_col150[139];
   data_col150[141] <= data_col150[140];
   data_col150[142] <= data_col150[141];
   data_col150[143] <= data_col150[142];
   data_col150[144] <= data_col150[143];
   data_col150[145] <= data_col150[144];
   data_col150[146] <= data_col150[145];
   data_col150[147] <= data_col150[146];
   data_col150[148] <= data_col150[147];
   data_col150[149] <= data_col150[148];
   data_col150[150] <= data_col150[149];

   data_col151[1] <= data[14];
   data_col151[2] <= data_col151[1];
   data_col151[3] <= data_col151[2];
   data_col151[4] <= data_col151[3];
   data_col151[5] <= data_col151[4];
   data_col151[6] <= data_col151[5];
   data_col151[7] <= data_col151[6];
   data_col151[8] <= data_col151[7];
   data_col151[9] <= data_col151[8];
   data_col151[10] <= data_col151[9];
   data_col151[11] <= data_col151[10];
   data_col151[12] <= data_col151[11];
   data_col151[13] <= data_col151[12];
   data_col151[14] <= data_col151[13];
   data_col151[15] <= data_col151[14];
   data_col151[16] <= data_col151[15];
   data_col151[17] <= data_col151[16];
   data_col151[18] <= data_col151[17];
   data_col151[19] <= data_col151[18];
   data_col151[20] <= data_col151[19];
   data_col151[21] <= data_col151[20];
   data_col151[22] <= data_col151[21];
   data_col151[23] <= data_col151[22];
   data_col151[24] <= data_col151[23];
   data_col151[25] <= data_col151[24];
   data_col151[26] <= data_col151[25];
   data_col151[27] <= data_col151[26];
   data_col151[28] <= data_col151[27];
   data_col151[29] <= data_col151[28];
   data_col151[30] <= data_col151[29];
   data_col151[31] <= data_col151[30];
   data_col151[32] <= data_col151[31];
   data_col151[33] <= data_col151[32];
   data_col151[34] <= data_col151[33];
   data_col151[35] <= data_col151[34];
   data_col151[36] <= data_col151[35];
   data_col151[37] <= data_col151[36];
   data_col151[38] <= data_col151[37];
   data_col151[39] <= data_col151[38];
   data_col151[40] <= data_col151[39];
   data_col151[41] <= data_col151[40];
   data_col151[42] <= data_col151[41];
   data_col151[43] <= data_col151[42];
   data_col151[44] <= data_col151[43];
   data_col151[45] <= data_col151[44];
   data_col151[46] <= data_col151[45];
   data_col151[47] <= data_col151[46];
   data_col151[48] <= data_col151[47];
   data_col151[49] <= data_col151[48];
   data_col151[50] <= data_col151[49];
   data_col151[51] <= data_col151[50];
   data_col151[52] <= data_col151[51];
   data_col151[53] <= data_col151[52];
   data_col151[54] <= data_col151[53];
   data_col151[55] <= data_col151[54];
   data_col151[56] <= data_col151[55];
   data_col151[57] <= data_col151[56];
   data_col151[58] <= data_col151[57];
   data_col151[59] <= data_col151[58];
   data_col151[60] <= data_col151[59];
   data_col151[61] <= data_col151[60];
   data_col151[62] <= data_col151[61];
   data_col151[63] <= data_col151[62];
   data_col151[64] <= data_col151[63];
   data_col151[65] <= data_col151[64];
   data_col151[66] <= data_col151[65];
   data_col151[67] <= data_col151[66];
   data_col151[68] <= data_col151[67];
   data_col151[69] <= data_col151[68];
   data_col151[70] <= data_col151[69];
   data_col151[71] <= data_col151[70];
   data_col151[72] <= data_col151[71];
   data_col151[73] <= data_col151[72];
   data_col151[74] <= data_col151[73];
   data_col151[75] <= data_col151[74];
   data_col151[76] <= data_col151[75];
   data_col151[77] <= data_col151[76];
   data_col151[78] <= data_col151[77];
   data_col151[79] <= data_col151[78];
   data_col151[80] <= data_col151[79];
   data_col151[81] <= data_col151[80];
   data_col151[82] <= data_col151[81];
   data_col151[83] <= data_col151[82];
   data_col151[84] <= data_col151[83];
   data_col151[85] <= data_col151[84];
   data_col151[86] <= data_col151[85];
   data_col151[87] <= data_col151[86];
   data_col151[88] <= data_col151[87];
   data_col151[89] <= data_col151[88];
   data_col151[90] <= data_col151[89];
   data_col151[91] <= data_col151[90];
   data_col151[92] <= data_col151[91];
   data_col151[93] <= data_col151[92];
   data_col151[94] <= data_col151[93];
   data_col151[95] <= data_col151[94];
   data_col151[96] <= data_col151[95];
   data_col151[97] <= data_col151[96];
   data_col151[98] <= data_col151[97];
   data_col151[99] <= data_col151[98];
   data_col151[100] <= data_col151[99];
   data_col151[101] <= data_col151[100];
   data_col151[102] <= data_col151[101];
   data_col151[103] <= data_col151[102];
   data_col151[104] <= data_col151[103];
   data_col151[105] <= data_col151[104];
   data_col151[106] <= data_col151[105];
   data_col151[107] <= data_col151[106];
   data_col151[108] <= data_col151[107];
   data_col151[109] <= data_col151[108];
   data_col151[110] <= data_col151[109];
   data_col151[111] <= data_col151[110];
   data_col151[112] <= data_col151[111];
   data_col151[113] <= data_col151[112];
   data_col151[114] <= data_col151[113];
   data_col151[115] <= data_col151[114];
   data_col151[116] <= data_col151[115];
   data_col151[117] <= data_col151[116];
   data_col151[118] <= data_col151[117];
   data_col151[119] <= data_col151[118];
   data_col151[120] <= data_col151[119];
   data_col151[121] <= data_col151[120];
   data_col151[122] <= data_col151[121];
   data_col151[123] <= data_col151[122];
   data_col151[124] <= data_col151[123];
   data_col151[125] <= data_col151[124];
   data_col151[126] <= data_col151[125];
   data_col151[127] <= data_col151[126];
   data_col151[128] <= data_col151[127];
   data_col151[129] <= data_col151[128];
   data_col151[130] <= data_col151[129];
   data_col151[131] <= data_col151[130];
   data_col151[132] <= data_col151[131];
   data_col151[133] <= data_col151[132];
   data_col151[134] <= data_col151[133];
   data_col151[135] <= data_col151[134];
   data_col151[136] <= data_col151[135];
   data_col151[137] <= data_col151[136];
   data_col151[138] <= data_col151[137];
   data_col151[139] <= data_col151[138];
   data_col151[140] <= data_col151[139];
   data_col151[141] <= data_col151[140];
   data_col151[142] <= data_col151[141];
   data_col151[143] <= data_col151[142];
   data_col151[144] <= data_col151[143];
   data_col151[145] <= data_col151[144];
   data_col151[146] <= data_col151[145];
   data_col151[147] <= data_col151[146];
   data_col151[148] <= data_col151[147];
   data_col151[149] <= data_col151[148];
   data_col151[150] <= data_col151[149];
   data_col151[151] <= data_col151[150];

   data_col152[1] <= data[13];
   data_col152[2] <= data_col152[1];
   data_col152[3] <= data_col152[2];
   data_col152[4] <= data_col152[3];
   data_col152[5] <= data_col152[4];
   data_col152[6] <= data_col152[5];
   data_col152[7] <= data_col152[6];
   data_col152[8] <= data_col152[7];
   data_col152[9] <= data_col152[8];
   data_col152[10] <= data_col152[9];
   data_col152[11] <= data_col152[10];
   data_col152[12] <= data_col152[11];
   data_col152[13] <= data_col152[12];
   data_col152[14] <= data_col152[13];
   data_col152[15] <= data_col152[14];
   data_col152[16] <= data_col152[15];
   data_col152[17] <= data_col152[16];
   data_col152[18] <= data_col152[17];
   data_col152[19] <= data_col152[18];
   data_col152[20] <= data_col152[19];
   data_col152[21] <= data_col152[20];
   data_col152[22] <= data_col152[21];
   data_col152[23] <= data_col152[22];
   data_col152[24] <= data_col152[23];
   data_col152[25] <= data_col152[24];
   data_col152[26] <= data_col152[25];
   data_col152[27] <= data_col152[26];
   data_col152[28] <= data_col152[27];
   data_col152[29] <= data_col152[28];
   data_col152[30] <= data_col152[29];
   data_col152[31] <= data_col152[30];
   data_col152[32] <= data_col152[31];
   data_col152[33] <= data_col152[32];
   data_col152[34] <= data_col152[33];
   data_col152[35] <= data_col152[34];
   data_col152[36] <= data_col152[35];
   data_col152[37] <= data_col152[36];
   data_col152[38] <= data_col152[37];
   data_col152[39] <= data_col152[38];
   data_col152[40] <= data_col152[39];
   data_col152[41] <= data_col152[40];
   data_col152[42] <= data_col152[41];
   data_col152[43] <= data_col152[42];
   data_col152[44] <= data_col152[43];
   data_col152[45] <= data_col152[44];
   data_col152[46] <= data_col152[45];
   data_col152[47] <= data_col152[46];
   data_col152[48] <= data_col152[47];
   data_col152[49] <= data_col152[48];
   data_col152[50] <= data_col152[49];
   data_col152[51] <= data_col152[50];
   data_col152[52] <= data_col152[51];
   data_col152[53] <= data_col152[52];
   data_col152[54] <= data_col152[53];
   data_col152[55] <= data_col152[54];
   data_col152[56] <= data_col152[55];
   data_col152[57] <= data_col152[56];
   data_col152[58] <= data_col152[57];
   data_col152[59] <= data_col152[58];
   data_col152[60] <= data_col152[59];
   data_col152[61] <= data_col152[60];
   data_col152[62] <= data_col152[61];
   data_col152[63] <= data_col152[62];
   data_col152[64] <= data_col152[63];
   data_col152[65] <= data_col152[64];
   data_col152[66] <= data_col152[65];
   data_col152[67] <= data_col152[66];
   data_col152[68] <= data_col152[67];
   data_col152[69] <= data_col152[68];
   data_col152[70] <= data_col152[69];
   data_col152[71] <= data_col152[70];
   data_col152[72] <= data_col152[71];
   data_col152[73] <= data_col152[72];
   data_col152[74] <= data_col152[73];
   data_col152[75] <= data_col152[74];
   data_col152[76] <= data_col152[75];
   data_col152[77] <= data_col152[76];
   data_col152[78] <= data_col152[77];
   data_col152[79] <= data_col152[78];
   data_col152[80] <= data_col152[79];
   data_col152[81] <= data_col152[80];
   data_col152[82] <= data_col152[81];
   data_col152[83] <= data_col152[82];
   data_col152[84] <= data_col152[83];
   data_col152[85] <= data_col152[84];
   data_col152[86] <= data_col152[85];
   data_col152[87] <= data_col152[86];
   data_col152[88] <= data_col152[87];
   data_col152[89] <= data_col152[88];
   data_col152[90] <= data_col152[89];
   data_col152[91] <= data_col152[90];
   data_col152[92] <= data_col152[91];
   data_col152[93] <= data_col152[92];
   data_col152[94] <= data_col152[93];
   data_col152[95] <= data_col152[94];
   data_col152[96] <= data_col152[95];
   data_col152[97] <= data_col152[96];
   data_col152[98] <= data_col152[97];
   data_col152[99] <= data_col152[98];
   data_col152[100] <= data_col152[99];
   data_col152[101] <= data_col152[100];
   data_col152[102] <= data_col152[101];
   data_col152[103] <= data_col152[102];
   data_col152[104] <= data_col152[103];
   data_col152[105] <= data_col152[104];
   data_col152[106] <= data_col152[105];
   data_col152[107] <= data_col152[106];
   data_col152[108] <= data_col152[107];
   data_col152[109] <= data_col152[108];
   data_col152[110] <= data_col152[109];
   data_col152[111] <= data_col152[110];
   data_col152[112] <= data_col152[111];
   data_col152[113] <= data_col152[112];
   data_col152[114] <= data_col152[113];
   data_col152[115] <= data_col152[114];
   data_col152[116] <= data_col152[115];
   data_col152[117] <= data_col152[116];
   data_col152[118] <= data_col152[117];
   data_col152[119] <= data_col152[118];
   data_col152[120] <= data_col152[119];
   data_col152[121] <= data_col152[120];
   data_col152[122] <= data_col152[121];
   data_col152[123] <= data_col152[122];
   data_col152[124] <= data_col152[123];
   data_col152[125] <= data_col152[124];
   data_col152[126] <= data_col152[125];
   data_col152[127] <= data_col152[126];
   data_col152[128] <= data_col152[127];
   data_col152[129] <= data_col152[128];
   data_col152[130] <= data_col152[129];
   data_col152[131] <= data_col152[130];
   data_col152[132] <= data_col152[131];
   data_col152[133] <= data_col152[132];
   data_col152[134] <= data_col152[133];
   data_col152[135] <= data_col152[134];
   data_col152[136] <= data_col152[135];
   data_col152[137] <= data_col152[136];
   data_col152[138] <= data_col152[137];
   data_col152[139] <= data_col152[138];
   data_col152[140] <= data_col152[139];
   data_col152[141] <= data_col152[140];
   data_col152[142] <= data_col152[141];
   data_col152[143] <= data_col152[142];
   data_col152[144] <= data_col152[143];
   data_col152[145] <= data_col152[144];
   data_col152[146] <= data_col152[145];
   data_col152[147] <= data_col152[146];
   data_col152[148] <= data_col152[147];
   data_col152[149] <= data_col152[148];
   data_col152[150] <= data_col152[149];
   data_col152[151] <= data_col152[150];
   data_col152[152] <= data_col152[151];

   data_col153[1] <= data[12];
   data_col153[2] <= data_col153[1];
   data_col153[3] <= data_col153[2];
   data_col153[4] <= data_col153[3];
   data_col153[5] <= data_col153[4];
   data_col153[6] <= data_col153[5];
   data_col153[7] <= data_col153[6];
   data_col153[8] <= data_col153[7];
   data_col153[9] <= data_col153[8];
   data_col153[10] <= data_col153[9];
   data_col153[11] <= data_col153[10];
   data_col153[12] <= data_col153[11];
   data_col153[13] <= data_col153[12];
   data_col153[14] <= data_col153[13];
   data_col153[15] <= data_col153[14];
   data_col153[16] <= data_col153[15];
   data_col153[17] <= data_col153[16];
   data_col153[18] <= data_col153[17];
   data_col153[19] <= data_col153[18];
   data_col153[20] <= data_col153[19];
   data_col153[21] <= data_col153[20];
   data_col153[22] <= data_col153[21];
   data_col153[23] <= data_col153[22];
   data_col153[24] <= data_col153[23];
   data_col153[25] <= data_col153[24];
   data_col153[26] <= data_col153[25];
   data_col153[27] <= data_col153[26];
   data_col153[28] <= data_col153[27];
   data_col153[29] <= data_col153[28];
   data_col153[30] <= data_col153[29];
   data_col153[31] <= data_col153[30];
   data_col153[32] <= data_col153[31];
   data_col153[33] <= data_col153[32];
   data_col153[34] <= data_col153[33];
   data_col153[35] <= data_col153[34];
   data_col153[36] <= data_col153[35];
   data_col153[37] <= data_col153[36];
   data_col153[38] <= data_col153[37];
   data_col153[39] <= data_col153[38];
   data_col153[40] <= data_col153[39];
   data_col153[41] <= data_col153[40];
   data_col153[42] <= data_col153[41];
   data_col153[43] <= data_col153[42];
   data_col153[44] <= data_col153[43];
   data_col153[45] <= data_col153[44];
   data_col153[46] <= data_col153[45];
   data_col153[47] <= data_col153[46];
   data_col153[48] <= data_col153[47];
   data_col153[49] <= data_col153[48];
   data_col153[50] <= data_col153[49];
   data_col153[51] <= data_col153[50];
   data_col153[52] <= data_col153[51];
   data_col153[53] <= data_col153[52];
   data_col153[54] <= data_col153[53];
   data_col153[55] <= data_col153[54];
   data_col153[56] <= data_col153[55];
   data_col153[57] <= data_col153[56];
   data_col153[58] <= data_col153[57];
   data_col153[59] <= data_col153[58];
   data_col153[60] <= data_col153[59];
   data_col153[61] <= data_col153[60];
   data_col153[62] <= data_col153[61];
   data_col153[63] <= data_col153[62];
   data_col153[64] <= data_col153[63];
   data_col153[65] <= data_col153[64];
   data_col153[66] <= data_col153[65];
   data_col153[67] <= data_col153[66];
   data_col153[68] <= data_col153[67];
   data_col153[69] <= data_col153[68];
   data_col153[70] <= data_col153[69];
   data_col153[71] <= data_col153[70];
   data_col153[72] <= data_col153[71];
   data_col153[73] <= data_col153[72];
   data_col153[74] <= data_col153[73];
   data_col153[75] <= data_col153[74];
   data_col153[76] <= data_col153[75];
   data_col153[77] <= data_col153[76];
   data_col153[78] <= data_col153[77];
   data_col153[79] <= data_col153[78];
   data_col153[80] <= data_col153[79];
   data_col153[81] <= data_col153[80];
   data_col153[82] <= data_col153[81];
   data_col153[83] <= data_col153[82];
   data_col153[84] <= data_col153[83];
   data_col153[85] <= data_col153[84];
   data_col153[86] <= data_col153[85];
   data_col153[87] <= data_col153[86];
   data_col153[88] <= data_col153[87];
   data_col153[89] <= data_col153[88];
   data_col153[90] <= data_col153[89];
   data_col153[91] <= data_col153[90];
   data_col153[92] <= data_col153[91];
   data_col153[93] <= data_col153[92];
   data_col153[94] <= data_col153[93];
   data_col153[95] <= data_col153[94];
   data_col153[96] <= data_col153[95];
   data_col153[97] <= data_col153[96];
   data_col153[98] <= data_col153[97];
   data_col153[99] <= data_col153[98];
   data_col153[100] <= data_col153[99];
   data_col153[101] <= data_col153[100];
   data_col153[102] <= data_col153[101];
   data_col153[103] <= data_col153[102];
   data_col153[104] <= data_col153[103];
   data_col153[105] <= data_col153[104];
   data_col153[106] <= data_col153[105];
   data_col153[107] <= data_col153[106];
   data_col153[108] <= data_col153[107];
   data_col153[109] <= data_col153[108];
   data_col153[110] <= data_col153[109];
   data_col153[111] <= data_col153[110];
   data_col153[112] <= data_col153[111];
   data_col153[113] <= data_col153[112];
   data_col153[114] <= data_col153[113];
   data_col153[115] <= data_col153[114];
   data_col153[116] <= data_col153[115];
   data_col153[117] <= data_col153[116];
   data_col153[118] <= data_col153[117];
   data_col153[119] <= data_col153[118];
   data_col153[120] <= data_col153[119];
   data_col153[121] <= data_col153[120];
   data_col153[122] <= data_col153[121];
   data_col153[123] <= data_col153[122];
   data_col153[124] <= data_col153[123];
   data_col153[125] <= data_col153[124];
   data_col153[126] <= data_col153[125];
   data_col153[127] <= data_col153[126];
   data_col153[128] <= data_col153[127];
   data_col153[129] <= data_col153[128];
   data_col153[130] <= data_col153[129];
   data_col153[131] <= data_col153[130];
   data_col153[132] <= data_col153[131];
   data_col153[133] <= data_col153[132];
   data_col153[134] <= data_col153[133];
   data_col153[135] <= data_col153[134];
   data_col153[136] <= data_col153[135];
   data_col153[137] <= data_col153[136];
   data_col153[138] <= data_col153[137];
   data_col153[139] <= data_col153[138];
   data_col153[140] <= data_col153[139];
   data_col153[141] <= data_col153[140];
   data_col153[142] <= data_col153[141];
   data_col153[143] <= data_col153[142];
   data_col153[144] <= data_col153[143];
   data_col153[145] <= data_col153[144];
   data_col153[146] <= data_col153[145];
   data_col153[147] <= data_col153[146];
   data_col153[148] <= data_col153[147];
   data_col153[149] <= data_col153[148];
   data_col153[150] <= data_col153[149];
   data_col153[151] <= data_col153[150];
   data_col153[152] <= data_col153[151];
   data_col153[153] <= data_col153[152];

   data_col154[1] <= data[11];
   data_col154[2] <= data_col154[1];
   data_col154[3] <= data_col154[2];
   data_col154[4] <= data_col154[3];
   data_col154[5] <= data_col154[4];
   data_col154[6] <= data_col154[5];
   data_col154[7] <= data_col154[6];
   data_col154[8] <= data_col154[7];
   data_col154[9] <= data_col154[8];
   data_col154[10] <= data_col154[9];
   data_col154[11] <= data_col154[10];
   data_col154[12] <= data_col154[11];
   data_col154[13] <= data_col154[12];
   data_col154[14] <= data_col154[13];
   data_col154[15] <= data_col154[14];
   data_col154[16] <= data_col154[15];
   data_col154[17] <= data_col154[16];
   data_col154[18] <= data_col154[17];
   data_col154[19] <= data_col154[18];
   data_col154[20] <= data_col154[19];
   data_col154[21] <= data_col154[20];
   data_col154[22] <= data_col154[21];
   data_col154[23] <= data_col154[22];
   data_col154[24] <= data_col154[23];
   data_col154[25] <= data_col154[24];
   data_col154[26] <= data_col154[25];
   data_col154[27] <= data_col154[26];
   data_col154[28] <= data_col154[27];
   data_col154[29] <= data_col154[28];
   data_col154[30] <= data_col154[29];
   data_col154[31] <= data_col154[30];
   data_col154[32] <= data_col154[31];
   data_col154[33] <= data_col154[32];
   data_col154[34] <= data_col154[33];
   data_col154[35] <= data_col154[34];
   data_col154[36] <= data_col154[35];
   data_col154[37] <= data_col154[36];
   data_col154[38] <= data_col154[37];
   data_col154[39] <= data_col154[38];
   data_col154[40] <= data_col154[39];
   data_col154[41] <= data_col154[40];
   data_col154[42] <= data_col154[41];
   data_col154[43] <= data_col154[42];
   data_col154[44] <= data_col154[43];
   data_col154[45] <= data_col154[44];
   data_col154[46] <= data_col154[45];
   data_col154[47] <= data_col154[46];
   data_col154[48] <= data_col154[47];
   data_col154[49] <= data_col154[48];
   data_col154[50] <= data_col154[49];
   data_col154[51] <= data_col154[50];
   data_col154[52] <= data_col154[51];
   data_col154[53] <= data_col154[52];
   data_col154[54] <= data_col154[53];
   data_col154[55] <= data_col154[54];
   data_col154[56] <= data_col154[55];
   data_col154[57] <= data_col154[56];
   data_col154[58] <= data_col154[57];
   data_col154[59] <= data_col154[58];
   data_col154[60] <= data_col154[59];
   data_col154[61] <= data_col154[60];
   data_col154[62] <= data_col154[61];
   data_col154[63] <= data_col154[62];
   data_col154[64] <= data_col154[63];
   data_col154[65] <= data_col154[64];
   data_col154[66] <= data_col154[65];
   data_col154[67] <= data_col154[66];
   data_col154[68] <= data_col154[67];
   data_col154[69] <= data_col154[68];
   data_col154[70] <= data_col154[69];
   data_col154[71] <= data_col154[70];
   data_col154[72] <= data_col154[71];
   data_col154[73] <= data_col154[72];
   data_col154[74] <= data_col154[73];
   data_col154[75] <= data_col154[74];
   data_col154[76] <= data_col154[75];
   data_col154[77] <= data_col154[76];
   data_col154[78] <= data_col154[77];
   data_col154[79] <= data_col154[78];
   data_col154[80] <= data_col154[79];
   data_col154[81] <= data_col154[80];
   data_col154[82] <= data_col154[81];
   data_col154[83] <= data_col154[82];
   data_col154[84] <= data_col154[83];
   data_col154[85] <= data_col154[84];
   data_col154[86] <= data_col154[85];
   data_col154[87] <= data_col154[86];
   data_col154[88] <= data_col154[87];
   data_col154[89] <= data_col154[88];
   data_col154[90] <= data_col154[89];
   data_col154[91] <= data_col154[90];
   data_col154[92] <= data_col154[91];
   data_col154[93] <= data_col154[92];
   data_col154[94] <= data_col154[93];
   data_col154[95] <= data_col154[94];
   data_col154[96] <= data_col154[95];
   data_col154[97] <= data_col154[96];
   data_col154[98] <= data_col154[97];
   data_col154[99] <= data_col154[98];
   data_col154[100] <= data_col154[99];
   data_col154[101] <= data_col154[100];
   data_col154[102] <= data_col154[101];
   data_col154[103] <= data_col154[102];
   data_col154[104] <= data_col154[103];
   data_col154[105] <= data_col154[104];
   data_col154[106] <= data_col154[105];
   data_col154[107] <= data_col154[106];
   data_col154[108] <= data_col154[107];
   data_col154[109] <= data_col154[108];
   data_col154[110] <= data_col154[109];
   data_col154[111] <= data_col154[110];
   data_col154[112] <= data_col154[111];
   data_col154[113] <= data_col154[112];
   data_col154[114] <= data_col154[113];
   data_col154[115] <= data_col154[114];
   data_col154[116] <= data_col154[115];
   data_col154[117] <= data_col154[116];
   data_col154[118] <= data_col154[117];
   data_col154[119] <= data_col154[118];
   data_col154[120] <= data_col154[119];
   data_col154[121] <= data_col154[120];
   data_col154[122] <= data_col154[121];
   data_col154[123] <= data_col154[122];
   data_col154[124] <= data_col154[123];
   data_col154[125] <= data_col154[124];
   data_col154[126] <= data_col154[125];
   data_col154[127] <= data_col154[126];
   data_col154[128] <= data_col154[127];
   data_col154[129] <= data_col154[128];
   data_col154[130] <= data_col154[129];
   data_col154[131] <= data_col154[130];
   data_col154[132] <= data_col154[131];
   data_col154[133] <= data_col154[132];
   data_col154[134] <= data_col154[133];
   data_col154[135] <= data_col154[134];
   data_col154[136] <= data_col154[135];
   data_col154[137] <= data_col154[136];
   data_col154[138] <= data_col154[137];
   data_col154[139] <= data_col154[138];
   data_col154[140] <= data_col154[139];
   data_col154[141] <= data_col154[140];
   data_col154[142] <= data_col154[141];
   data_col154[143] <= data_col154[142];
   data_col154[144] <= data_col154[143];
   data_col154[145] <= data_col154[144];
   data_col154[146] <= data_col154[145];
   data_col154[147] <= data_col154[146];
   data_col154[148] <= data_col154[147];
   data_col154[149] <= data_col154[148];
   data_col154[150] <= data_col154[149];
   data_col154[151] <= data_col154[150];
   data_col154[152] <= data_col154[151];
   data_col154[153] <= data_col154[152];
   data_col154[154] <= data_col154[153];

   data_col155[1] <= data[10];
   data_col155[2] <= data_col155[1];
   data_col155[3] <= data_col155[2];
   data_col155[4] <= data_col155[3];
   data_col155[5] <= data_col155[4];
   data_col155[6] <= data_col155[5];
   data_col155[7] <= data_col155[6];
   data_col155[8] <= data_col155[7];
   data_col155[9] <= data_col155[8];
   data_col155[10] <= data_col155[9];
   data_col155[11] <= data_col155[10];
   data_col155[12] <= data_col155[11];
   data_col155[13] <= data_col155[12];
   data_col155[14] <= data_col155[13];
   data_col155[15] <= data_col155[14];
   data_col155[16] <= data_col155[15];
   data_col155[17] <= data_col155[16];
   data_col155[18] <= data_col155[17];
   data_col155[19] <= data_col155[18];
   data_col155[20] <= data_col155[19];
   data_col155[21] <= data_col155[20];
   data_col155[22] <= data_col155[21];
   data_col155[23] <= data_col155[22];
   data_col155[24] <= data_col155[23];
   data_col155[25] <= data_col155[24];
   data_col155[26] <= data_col155[25];
   data_col155[27] <= data_col155[26];
   data_col155[28] <= data_col155[27];
   data_col155[29] <= data_col155[28];
   data_col155[30] <= data_col155[29];
   data_col155[31] <= data_col155[30];
   data_col155[32] <= data_col155[31];
   data_col155[33] <= data_col155[32];
   data_col155[34] <= data_col155[33];
   data_col155[35] <= data_col155[34];
   data_col155[36] <= data_col155[35];
   data_col155[37] <= data_col155[36];
   data_col155[38] <= data_col155[37];
   data_col155[39] <= data_col155[38];
   data_col155[40] <= data_col155[39];
   data_col155[41] <= data_col155[40];
   data_col155[42] <= data_col155[41];
   data_col155[43] <= data_col155[42];
   data_col155[44] <= data_col155[43];
   data_col155[45] <= data_col155[44];
   data_col155[46] <= data_col155[45];
   data_col155[47] <= data_col155[46];
   data_col155[48] <= data_col155[47];
   data_col155[49] <= data_col155[48];
   data_col155[50] <= data_col155[49];
   data_col155[51] <= data_col155[50];
   data_col155[52] <= data_col155[51];
   data_col155[53] <= data_col155[52];
   data_col155[54] <= data_col155[53];
   data_col155[55] <= data_col155[54];
   data_col155[56] <= data_col155[55];
   data_col155[57] <= data_col155[56];
   data_col155[58] <= data_col155[57];
   data_col155[59] <= data_col155[58];
   data_col155[60] <= data_col155[59];
   data_col155[61] <= data_col155[60];
   data_col155[62] <= data_col155[61];
   data_col155[63] <= data_col155[62];
   data_col155[64] <= data_col155[63];
   data_col155[65] <= data_col155[64];
   data_col155[66] <= data_col155[65];
   data_col155[67] <= data_col155[66];
   data_col155[68] <= data_col155[67];
   data_col155[69] <= data_col155[68];
   data_col155[70] <= data_col155[69];
   data_col155[71] <= data_col155[70];
   data_col155[72] <= data_col155[71];
   data_col155[73] <= data_col155[72];
   data_col155[74] <= data_col155[73];
   data_col155[75] <= data_col155[74];
   data_col155[76] <= data_col155[75];
   data_col155[77] <= data_col155[76];
   data_col155[78] <= data_col155[77];
   data_col155[79] <= data_col155[78];
   data_col155[80] <= data_col155[79];
   data_col155[81] <= data_col155[80];
   data_col155[82] <= data_col155[81];
   data_col155[83] <= data_col155[82];
   data_col155[84] <= data_col155[83];
   data_col155[85] <= data_col155[84];
   data_col155[86] <= data_col155[85];
   data_col155[87] <= data_col155[86];
   data_col155[88] <= data_col155[87];
   data_col155[89] <= data_col155[88];
   data_col155[90] <= data_col155[89];
   data_col155[91] <= data_col155[90];
   data_col155[92] <= data_col155[91];
   data_col155[93] <= data_col155[92];
   data_col155[94] <= data_col155[93];
   data_col155[95] <= data_col155[94];
   data_col155[96] <= data_col155[95];
   data_col155[97] <= data_col155[96];
   data_col155[98] <= data_col155[97];
   data_col155[99] <= data_col155[98];
   data_col155[100] <= data_col155[99];
   data_col155[101] <= data_col155[100];
   data_col155[102] <= data_col155[101];
   data_col155[103] <= data_col155[102];
   data_col155[104] <= data_col155[103];
   data_col155[105] <= data_col155[104];
   data_col155[106] <= data_col155[105];
   data_col155[107] <= data_col155[106];
   data_col155[108] <= data_col155[107];
   data_col155[109] <= data_col155[108];
   data_col155[110] <= data_col155[109];
   data_col155[111] <= data_col155[110];
   data_col155[112] <= data_col155[111];
   data_col155[113] <= data_col155[112];
   data_col155[114] <= data_col155[113];
   data_col155[115] <= data_col155[114];
   data_col155[116] <= data_col155[115];
   data_col155[117] <= data_col155[116];
   data_col155[118] <= data_col155[117];
   data_col155[119] <= data_col155[118];
   data_col155[120] <= data_col155[119];
   data_col155[121] <= data_col155[120];
   data_col155[122] <= data_col155[121];
   data_col155[123] <= data_col155[122];
   data_col155[124] <= data_col155[123];
   data_col155[125] <= data_col155[124];
   data_col155[126] <= data_col155[125];
   data_col155[127] <= data_col155[126];
   data_col155[128] <= data_col155[127];
   data_col155[129] <= data_col155[128];
   data_col155[130] <= data_col155[129];
   data_col155[131] <= data_col155[130];
   data_col155[132] <= data_col155[131];
   data_col155[133] <= data_col155[132];
   data_col155[134] <= data_col155[133];
   data_col155[135] <= data_col155[134];
   data_col155[136] <= data_col155[135];
   data_col155[137] <= data_col155[136];
   data_col155[138] <= data_col155[137];
   data_col155[139] <= data_col155[138];
   data_col155[140] <= data_col155[139];
   data_col155[141] <= data_col155[140];
   data_col155[142] <= data_col155[141];
   data_col155[143] <= data_col155[142];
   data_col155[144] <= data_col155[143];
   data_col155[145] <= data_col155[144];
   data_col155[146] <= data_col155[145];
   data_col155[147] <= data_col155[146];
   data_col155[148] <= data_col155[147];
   data_col155[149] <= data_col155[148];
   data_col155[150] <= data_col155[149];
   data_col155[151] <= data_col155[150];
   data_col155[152] <= data_col155[151];
   data_col155[153] <= data_col155[152];
   data_col155[154] <= data_col155[153];
   data_col155[155] <= data_col155[154];

   data_col156[1] <= data[9];
   data_col156[2] <= data_col156[1];
   data_col156[3] <= data_col156[2];
   data_col156[4] <= data_col156[3];
   data_col156[5] <= data_col156[4];
   data_col156[6] <= data_col156[5];
   data_col156[7] <= data_col156[6];
   data_col156[8] <= data_col156[7];
   data_col156[9] <= data_col156[8];
   data_col156[10] <= data_col156[9];
   data_col156[11] <= data_col156[10];
   data_col156[12] <= data_col156[11];
   data_col156[13] <= data_col156[12];
   data_col156[14] <= data_col156[13];
   data_col156[15] <= data_col156[14];
   data_col156[16] <= data_col156[15];
   data_col156[17] <= data_col156[16];
   data_col156[18] <= data_col156[17];
   data_col156[19] <= data_col156[18];
   data_col156[20] <= data_col156[19];
   data_col156[21] <= data_col156[20];
   data_col156[22] <= data_col156[21];
   data_col156[23] <= data_col156[22];
   data_col156[24] <= data_col156[23];
   data_col156[25] <= data_col156[24];
   data_col156[26] <= data_col156[25];
   data_col156[27] <= data_col156[26];
   data_col156[28] <= data_col156[27];
   data_col156[29] <= data_col156[28];
   data_col156[30] <= data_col156[29];
   data_col156[31] <= data_col156[30];
   data_col156[32] <= data_col156[31];
   data_col156[33] <= data_col156[32];
   data_col156[34] <= data_col156[33];
   data_col156[35] <= data_col156[34];
   data_col156[36] <= data_col156[35];
   data_col156[37] <= data_col156[36];
   data_col156[38] <= data_col156[37];
   data_col156[39] <= data_col156[38];
   data_col156[40] <= data_col156[39];
   data_col156[41] <= data_col156[40];
   data_col156[42] <= data_col156[41];
   data_col156[43] <= data_col156[42];
   data_col156[44] <= data_col156[43];
   data_col156[45] <= data_col156[44];
   data_col156[46] <= data_col156[45];
   data_col156[47] <= data_col156[46];
   data_col156[48] <= data_col156[47];
   data_col156[49] <= data_col156[48];
   data_col156[50] <= data_col156[49];
   data_col156[51] <= data_col156[50];
   data_col156[52] <= data_col156[51];
   data_col156[53] <= data_col156[52];
   data_col156[54] <= data_col156[53];
   data_col156[55] <= data_col156[54];
   data_col156[56] <= data_col156[55];
   data_col156[57] <= data_col156[56];
   data_col156[58] <= data_col156[57];
   data_col156[59] <= data_col156[58];
   data_col156[60] <= data_col156[59];
   data_col156[61] <= data_col156[60];
   data_col156[62] <= data_col156[61];
   data_col156[63] <= data_col156[62];
   data_col156[64] <= data_col156[63];
   data_col156[65] <= data_col156[64];
   data_col156[66] <= data_col156[65];
   data_col156[67] <= data_col156[66];
   data_col156[68] <= data_col156[67];
   data_col156[69] <= data_col156[68];
   data_col156[70] <= data_col156[69];
   data_col156[71] <= data_col156[70];
   data_col156[72] <= data_col156[71];
   data_col156[73] <= data_col156[72];
   data_col156[74] <= data_col156[73];
   data_col156[75] <= data_col156[74];
   data_col156[76] <= data_col156[75];
   data_col156[77] <= data_col156[76];
   data_col156[78] <= data_col156[77];
   data_col156[79] <= data_col156[78];
   data_col156[80] <= data_col156[79];
   data_col156[81] <= data_col156[80];
   data_col156[82] <= data_col156[81];
   data_col156[83] <= data_col156[82];
   data_col156[84] <= data_col156[83];
   data_col156[85] <= data_col156[84];
   data_col156[86] <= data_col156[85];
   data_col156[87] <= data_col156[86];
   data_col156[88] <= data_col156[87];
   data_col156[89] <= data_col156[88];
   data_col156[90] <= data_col156[89];
   data_col156[91] <= data_col156[90];
   data_col156[92] <= data_col156[91];
   data_col156[93] <= data_col156[92];
   data_col156[94] <= data_col156[93];
   data_col156[95] <= data_col156[94];
   data_col156[96] <= data_col156[95];
   data_col156[97] <= data_col156[96];
   data_col156[98] <= data_col156[97];
   data_col156[99] <= data_col156[98];
   data_col156[100] <= data_col156[99];
   data_col156[101] <= data_col156[100];
   data_col156[102] <= data_col156[101];
   data_col156[103] <= data_col156[102];
   data_col156[104] <= data_col156[103];
   data_col156[105] <= data_col156[104];
   data_col156[106] <= data_col156[105];
   data_col156[107] <= data_col156[106];
   data_col156[108] <= data_col156[107];
   data_col156[109] <= data_col156[108];
   data_col156[110] <= data_col156[109];
   data_col156[111] <= data_col156[110];
   data_col156[112] <= data_col156[111];
   data_col156[113] <= data_col156[112];
   data_col156[114] <= data_col156[113];
   data_col156[115] <= data_col156[114];
   data_col156[116] <= data_col156[115];
   data_col156[117] <= data_col156[116];
   data_col156[118] <= data_col156[117];
   data_col156[119] <= data_col156[118];
   data_col156[120] <= data_col156[119];
   data_col156[121] <= data_col156[120];
   data_col156[122] <= data_col156[121];
   data_col156[123] <= data_col156[122];
   data_col156[124] <= data_col156[123];
   data_col156[125] <= data_col156[124];
   data_col156[126] <= data_col156[125];
   data_col156[127] <= data_col156[126];
   data_col156[128] <= data_col156[127];
   data_col156[129] <= data_col156[128];
   data_col156[130] <= data_col156[129];
   data_col156[131] <= data_col156[130];
   data_col156[132] <= data_col156[131];
   data_col156[133] <= data_col156[132];
   data_col156[134] <= data_col156[133];
   data_col156[135] <= data_col156[134];
   data_col156[136] <= data_col156[135];
   data_col156[137] <= data_col156[136];
   data_col156[138] <= data_col156[137];
   data_col156[139] <= data_col156[138];
   data_col156[140] <= data_col156[139];
   data_col156[141] <= data_col156[140];
   data_col156[142] <= data_col156[141];
   data_col156[143] <= data_col156[142];
   data_col156[144] <= data_col156[143];
   data_col156[145] <= data_col156[144];
   data_col156[146] <= data_col156[145];
   data_col156[147] <= data_col156[146];
   data_col156[148] <= data_col156[147];
   data_col156[149] <= data_col156[148];
   data_col156[150] <= data_col156[149];
   data_col156[151] <= data_col156[150];
   data_col156[152] <= data_col156[151];
   data_col156[153] <= data_col156[152];
   data_col156[154] <= data_col156[153];
   data_col156[155] <= data_col156[154];
   data_col156[156] <= data_col156[155];

   data_col157[1] <= data[8];
   data_col157[2] <= data_col157[1];
   data_col157[3] <= data_col157[2];
   data_col157[4] <= data_col157[3];
   data_col157[5] <= data_col157[4];
   data_col157[6] <= data_col157[5];
   data_col157[7] <= data_col157[6];
   data_col157[8] <= data_col157[7];
   data_col157[9] <= data_col157[8];
   data_col157[10] <= data_col157[9];
   data_col157[11] <= data_col157[10];
   data_col157[12] <= data_col157[11];
   data_col157[13] <= data_col157[12];
   data_col157[14] <= data_col157[13];
   data_col157[15] <= data_col157[14];
   data_col157[16] <= data_col157[15];
   data_col157[17] <= data_col157[16];
   data_col157[18] <= data_col157[17];
   data_col157[19] <= data_col157[18];
   data_col157[20] <= data_col157[19];
   data_col157[21] <= data_col157[20];
   data_col157[22] <= data_col157[21];
   data_col157[23] <= data_col157[22];
   data_col157[24] <= data_col157[23];
   data_col157[25] <= data_col157[24];
   data_col157[26] <= data_col157[25];
   data_col157[27] <= data_col157[26];
   data_col157[28] <= data_col157[27];
   data_col157[29] <= data_col157[28];
   data_col157[30] <= data_col157[29];
   data_col157[31] <= data_col157[30];
   data_col157[32] <= data_col157[31];
   data_col157[33] <= data_col157[32];
   data_col157[34] <= data_col157[33];
   data_col157[35] <= data_col157[34];
   data_col157[36] <= data_col157[35];
   data_col157[37] <= data_col157[36];
   data_col157[38] <= data_col157[37];
   data_col157[39] <= data_col157[38];
   data_col157[40] <= data_col157[39];
   data_col157[41] <= data_col157[40];
   data_col157[42] <= data_col157[41];
   data_col157[43] <= data_col157[42];
   data_col157[44] <= data_col157[43];
   data_col157[45] <= data_col157[44];
   data_col157[46] <= data_col157[45];
   data_col157[47] <= data_col157[46];
   data_col157[48] <= data_col157[47];
   data_col157[49] <= data_col157[48];
   data_col157[50] <= data_col157[49];
   data_col157[51] <= data_col157[50];
   data_col157[52] <= data_col157[51];
   data_col157[53] <= data_col157[52];
   data_col157[54] <= data_col157[53];
   data_col157[55] <= data_col157[54];
   data_col157[56] <= data_col157[55];
   data_col157[57] <= data_col157[56];
   data_col157[58] <= data_col157[57];
   data_col157[59] <= data_col157[58];
   data_col157[60] <= data_col157[59];
   data_col157[61] <= data_col157[60];
   data_col157[62] <= data_col157[61];
   data_col157[63] <= data_col157[62];
   data_col157[64] <= data_col157[63];
   data_col157[65] <= data_col157[64];
   data_col157[66] <= data_col157[65];
   data_col157[67] <= data_col157[66];
   data_col157[68] <= data_col157[67];
   data_col157[69] <= data_col157[68];
   data_col157[70] <= data_col157[69];
   data_col157[71] <= data_col157[70];
   data_col157[72] <= data_col157[71];
   data_col157[73] <= data_col157[72];
   data_col157[74] <= data_col157[73];
   data_col157[75] <= data_col157[74];
   data_col157[76] <= data_col157[75];
   data_col157[77] <= data_col157[76];
   data_col157[78] <= data_col157[77];
   data_col157[79] <= data_col157[78];
   data_col157[80] <= data_col157[79];
   data_col157[81] <= data_col157[80];
   data_col157[82] <= data_col157[81];
   data_col157[83] <= data_col157[82];
   data_col157[84] <= data_col157[83];
   data_col157[85] <= data_col157[84];
   data_col157[86] <= data_col157[85];
   data_col157[87] <= data_col157[86];
   data_col157[88] <= data_col157[87];
   data_col157[89] <= data_col157[88];
   data_col157[90] <= data_col157[89];
   data_col157[91] <= data_col157[90];
   data_col157[92] <= data_col157[91];
   data_col157[93] <= data_col157[92];
   data_col157[94] <= data_col157[93];
   data_col157[95] <= data_col157[94];
   data_col157[96] <= data_col157[95];
   data_col157[97] <= data_col157[96];
   data_col157[98] <= data_col157[97];
   data_col157[99] <= data_col157[98];
   data_col157[100] <= data_col157[99];
   data_col157[101] <= data_col157[100];
   data_col157[102] <= data_col157[101];
   data_col157[103] <= data_col157[102];
   data_col157[104] <= data_col157[103];
   data_col157[105] <= data_col157[104];
   data_col157[106] <= data_col157[105];
   data_col157[107] <= data_col157[106];
   data_col157[108] <= data_col157[107];
   data_col157[109] <= data_col157[108];
   data_col157[110] <= data_col157[109];
   data_col157[111] <= data_col157[110];
   data_col157[112] <= data_col157[111];
   data_col157[113] <= data_col157[112];
   data_col157[114] <= data_col157[113];
   data_col157[115] <= data_col157[114];
   data_col157[116] <= data_col157[115];
   data_col157[117] <= data_col157[116];
   data_col157[118] <= data_col157[117];
   data_col157[119] <= data_col157[118];
   data_col157[120] <= data_col157[119];
   data_col157[121] <= data_col157[120];
   data_col157[122] <= data_col157[121];
   data_col157[123] <= data_col157[122];
   data_col157[124] <= data_col157[123];
   data_col157[125] <= data_col157[124];
   data_col157[126] <= data_col157[125];
   data_col157[127] <= data_col157[126];
   data_col157[128] <= data_col157[127];
   data_col157[129] <= data_col157[128];
   data_col157[130] <= data_col157[129];
   data_col157[131] <= data_col157[130];
   data_col157[132] <= data_col157[131];
   data_col157[133] <= data_col157[132];
   data_col157[134] <= data_col157[133];
   data_col157[135] <= data_col157[134];
   data_col157[136] <= data_col157[135];
   data_col157[137] <= data_col157[136];
   data_col157[138] <= data_col157[137];
   data_col157[139] <= data_col157[138];
   data_col157[140] <= data_col157[139];
   data_col157[141] <= data_col157[140];
   data_col157[142] <= data_col157[141];
   data_col157[143] <= data_col157[142];
   data_col157[144] <= data_col157[143];
   data_col157[145] <= data_col157[144];
   data_col157[146] <= data_col157[145];
   data_col157[147] <= data_col157[146];
   data_col157[148] <= data_col157[147];
   data_col157[149] <= data_col157[148];
   data_col157[150] <= data_col157[149];
   data_col157[151] <= data_col157[150];
   data_col157[152] <= data_col157[151];
   data_col157[153] <= data_col157[152];
   data_col157[154] <= data_col157[153];
   data_col157[155] <= data_col157[154];
   data_col157[156] <= data_col157[155];
   data_col157[157] <= data_col157[156];

   data_col158[1] <= data[7];
   data_col158[2] <= data_col158[1];
   data_col158[3] <= data_col158[2];
   data_col158[4] <= data_col158[3];
   data_col158[5] <= data_col158[4];
   data_col158[6] <= data_col158[5];
   data_col158[7] <= data_col158[6];
   data_col158[8] <= data_col158[7];
   data_col158[9] <= data_col158[8];
   data_col158[10] <= data_col158[9];
   data_col158[11] <= data_col158[10];
   data_col158[12] <= data_col158[11];
   data_col158[13] <= data_col158[12];
   data_col158[14] <= data_col158[13];
   data_col158[15] <= data_col158[14];
   data_col158[16] <= data_col158[15];
   data_col158[17] <= data_col158[16];
   data_col158[18] <= data_col158[17];
   data_col158[19] <= data_col158[18];
   data_col158[20] <= data_col158[19];
   data_col158[21] <= data_col158[20];
   data_col158[22] <= data_col158[21];
   data_col158[23] <= data_col158[22];
   data_col158[24] <= data_col158[23];
   data_col158[25] <= data_col158[24];
   data_col158[26] <= data_col158[25];
   data_col158[27] <= data_col158[26];
   data_col158[28] <= data_col158[27];
   data_col158[29] <= data_col158[28];
   data_col158[30] <= data_col158[29];
   data_col158[31] <= data_col158[30];
   data_col158[32] <= data_col158[31];
   data_col158[33] <= data_col158[32];
   data_col158[34] <= data_col158[33];
   data_col158[35] <= data_col158[34];
   data_col158[36] <= data_col158[35];
   data_col158[37] <= data_col158[36];
   data_col158[38] <= data_col158[37];
   data_col158[39] <= data_col158[38];
   data_col158[40] <= data_col158[39];
   data_col158[41] <= data_col158[40];
   data_col158[42] <= data_col158[41];
   data_col158[43] <= data_col158[42];
   data_col158[44] <= data_col158[43];
   data_col158[45] <= data_col158[44];
   data_col158[46] <= data_col158[45];
   data_col158[47] <= data_col158[46];
   data_col158[48] <= data_col158[47];
   data_col158[49] <= data_col158[48];
   data_col158[50] <= data_col158[49];
   data_col158[51] <= data_col158[50];
   data_col158[52] <= data_col158[51];
   data_col158[53] <= data_col158[52];
   data_col158[54] <= data_col158[53];
   data_col158[55] <= data_col158[54];
   data_col158[56] <= data_col158[55];
   data_col158[57] <= data_col158[56];
   data_col158[58] <= data_col158[57];
   data_col158[59] <= data_col158[58];
   data_col158[60] <= data_col158[59];
   data_col158[61] <= data_col158[60];
   data_col158[62] <= data_col158[61];
   data_col158[63] <= data_col158[62];
   data_col158[64] <= data_col158[63];
   data_col158[65] <= data_col158[64];
   data_col158[66] <= data_col158[65];
   data_col158[67] <= data_col158[66];
   data_col158[68] <= data_col158[67];
   data_col158[69] <= data_col158[68];
   data_col158[70] <= data_col158[69];
   data_col158[71] <= data_col158[70];
   data_col158[72] <= data_col158[71];
   data_col158[73] <= data_col158[72];
   data_col158[74] <= data_col158[73];
   data_col158[75] <= data_col158[74];
   data_col158[76] <= data_col158[75];
   data_col158[77] <= data_col158[76];
   data_col158[78] <= data_col158[77];
   data_col158[79] <= data_col158[78];
   data_col158[80] <= data_col158[79];
   data_col158[81] <= data_col158[80];
   data_col158[82] <= data_col158[81];
   data_col158[83] <= data_col158[82];
   data_col158[84] <= data_col158[83];
   data_col158[85] <= data_col158[84];
   data_col158[86] <= data_col158[85];
   data_col158[87] <= data_col158[86];
   data_col158[88] <= data_col158[87];
   data_col158[89] <= data_col158[88];
   data_col158[90] <= data_col158[89];
   data_col158[91] <= data_col158[90];
   data_col158[92] <= data_col158[91];
   data_col158[93] <= data_col158[92];
   data_col158[94] <= data_col158[93];
   data_col158[95] <= data_col158[94];
   data_col158[96] <= data_col158[95];
   data_col158[97] <= data_col158[96];
   data_col158[98] <= data_col158[97];
   data_col158[99] <= data_col158[98];
   data_col158[100] <= data_col158[99];
   data_col158[101] <= data_col158[100];
   data_col158[102] <= data_col158[101];
   data_col158[103] <= data_col158[102];
   data_col158[104] <= data_col158[103];
   data_col158[105] <= data_col158[104];
   data_col158[106] <= data_col158[105];
   data_col158[107] <= data_col158[106];
   data_col158[108] <= data_col158[107];
   data_col158[109] <= data_col158[108];
   data_col158[110] <= data_col158[109];
   data_col158[111] <= data_col158[110];
   data_col158[112] <= data_col158[111];
   data_col158[113] <= data_col158[112];
   data_col158[114] <= data_col158[113];
   data_col158[115] <= data_col158[114];
   data_col158[116] <= data_col158[115];
   data_col158[117] <= data_col158[116];
   data_col158[118] <= data_col158[117];
   data_col158[119] <= data_col158[118];
   data_col158[120] <= data_col158[119];
   data_col158[121] <= data_col158[120];
   data_col158[122] <= data_col158[121];
   data_col158[123] <= data_col158[122];
   data_col158[124] <= data_col158[123];
   data_col158[125] <= data_col158[124];
   data_col158[126] <= data_col158[125];
   data_col158[127] <= data_col158[126];
   data_col158[128] <= data_col158[127];
   data_col158[129] <= data_col158[128];
   data_col158[130] <= data_col158[129];
   data_col158[131] <= data_col158[130];
   data_col158[132] <= data_col158[131];
   data_col158[133] <= data_col158[132];
   data_col158[134] <= data_col158[133];
   data_col158[135] <= data_col158[134];
   data_col158[136] <= data_col158[135];
   data_col158[137] <= data_col158[136];
   data_col158[138] <= data_col158[137];
   data_col158[139] <= data_col158[138];
   data_col158[140] <= data_col158[139];
   data_col158[141] <= data_col158[140];
   data_col158[142] <= data_col158[141];
   data_col158[143] <= data_col158[142];
   data_col158[144] <= data_col158[143];
   data_col158[145] <= data_col158[144];
   data_col158[146] <= data_col158[145];
   data_col158[147] <= data_col158[146];
   data_col158[148] <= data_col158[147];
   data_col158[149] <= data_col158[148];
   data_col158[150] <= data_col158[149];
   data_col158[151] <= data_col158[150];
   data_col158[152] <= data_col158[151];
   data_col158[153] <= data_col158[152];
   data_col158[154] <= data_col158[153];
   data_col158[155] <= data_col158[154];
   data_col158[156] <= data_col158[155];
   data_col158[157] <= data_col158[156];
   data_col158[158] <= data_col158[157];

   data_col159[1] <= data[6];
   data_col159[2] <= data_col159[1];
   data_col159[3] <= data_col159[2];
   data_col159[4] <= data_col159[3];
   data_col159[5] <= data_col159[4];
   data_col159[6] <= data_col159[5];
   data_col159[7] <= data_col159[6];
   data_col159[8] <= data_col159[7];
   data_col159[9] <= data_col159[8];
   data_col159[10] <= data_col159[9];
   data_col159[11] <= data_col159[10];
   data_col159[12] <= data_col159[11];
   data_col159[13] <= data_col159[12];
   data_col159[14] <= data_col159[13];
   data_col159[15] <= data_col159[14];
   data_col159[16] <= data_col159[15];
   data_col159[17] <= data_col159[16];
   data_col159[18] <= data_col159[17];
   data_col159[19] <= data_col159[18];
   data_col159[20] <= data_col159[19];
   data_col159[21] <= data_col159[20];
   data_col159[22] <= data_col159[21];
   data_col159[23] <= data_col159[22];
   data_col159[24] <= data_col159[23];
   data_col159[25] <= data_col159[24];
   data_col159[26] <= data_col159[25];
   data_col159[27] <= data_col159[26];
   data_col159[28] <= data_col159[27];
   data_col159[29] <= data_col159[28];
   data_col159[30] <= data_col159[29];
   data_col159[31] <= data_col159[30];
   data_col159[32] <= data_col159[31];
   data_col159[33] <= data_col159[32];
   data_col159[34] <= data_col159[33];
   data_col159[35] <= data_col159[34];
   data_col159[36] <= data_col159[35];
   data_col159[37] <= data_col159[36];
   data_col159[38] <= data_col159[37];
   data_col159[39] <= data_col159[38];
   data_col159[40] <= data_col159[39];
   data_col159[41] <= data_col159[40];
   data_col159[42] <= data_col159[41];
   data_col159[43] <= data_col159[42];
   data_col159[44] <= data_col159[43];
   data_col159[45] <= data_col159[44];
   data_col159[46] <= data_col159[45];
   data_col159[47] <= data_col159[46];
   data_col159[48] <= data_col159[47];
   data_col159[49] <= data_col159[48];
   data_col159[50] <= data_col159[49];
   data_col159[51] <= data_col159[50];
   data_col159[52] <= data_col159[51];
   data_col159[53] <= data_col159[52];
   data_col159[54] <= data_col159[53];
   data_col159[55] <= data_col159[54];
   data_col159[56] <= data_col159[55];
   data_col159[57] <= data_col159[56];
   data_col159[58] <= data_col159[57];
   data_col159[59] <= data_col159[58];
   data_col159[60] <= data_col159[59];
   data_col159[61] <= data_col159[60];
   data_col159[62] <= data_col159[61];
   data_col159[63] <= data_col159[62];
   data_col159[64] <= data_col159[63];
   data_col159[65] <= data_col159[64];
   data_col159[66] <= data_col159[65];
   data_col159[67] <= data_col159[66];
   data_col159[68] <= data_col159[67];
   data_col159[69] <= data_col159[68];
   data_col159[70] <= data_col159[69];
   data_col159[71] <= data_col159[70];
   data_col159[72] <= data_col159[71];
   data_col159[73] <= data_col159[72];
   data_col159[74] <= data_col159[73];
   data_col159[75] <= data_col159[74];
   data_col159[76] <= data_col159[75];
   data_col159[77] <= data_col159[76];
   data_col159[78] <= data_col159[77];
   data_col159[79] <= data_col159[78];
   data_col159[80] <= data_col159[79];
   data_col159[81] <= data_col159[80];
   data_col159[82] <= data_col159[81];
   data_col159[83] <= data_col159[82];
   data_col159[84] <= data_col159[83];
   data_col159[85] <= data_col159[84];
   data_col159[86] <= data_col159[85];
   data_col159[87] <= data_col159[86];
   data_col159[88] <= data_col159[87];
   data_col159[89] <= data_col159[88];
   data_col159[90] <= data_col159[89];
   data_col159[91] <= data_col159[90];
   data_col159[92] <= data_col159[91];
   data_col159[93] <= data_col159[92];
   data_col159[94] <= data_col159[93];
   data_col159[95] <= data_col159[94];
   data_col159[96] <= data_col159[95];
   data_col159[97] <= data_col159[96];
   data_col159[98] <= data_col159[97];
   data_col159[99] <= data_col159[98];
   data_col159[100] <= data_col159[99];
   data_col159[101] <= data_col159[100];
   data_col159[102] <= data_col159[101];
   data_col159[103] <= data_col159[102];
   data_col159[104] <= data_col159[103];
   data_col159[105] <= data_col159[104];
   data_col159[106] <= data_col159[105];
   data_col159[107] <= data_col159[106];
   data_col159[108] <= data_col159[107];
   data_col159[109] <= data_col159[108];
   data_col159[110] <= data_col159[109];
   data_col159[111] <= data_col159[110];
   data_col159[112] <= data_col159[111];
   data_col159[113] <= data_col159[112];
   data_col159[114] <= data_col159[113];
   data_col159[115] <= data_col159[114];
   data_col159[116] <= data_col159[115];
   data_col159[117] <= data_col159[116];
   data_col159[118] <= data_col159[117];
   data_col159[119] <= data_col159[118];
   data_col159[120] <= data_col159[119];
   data_col159[121] <= data_col159[120];
   data_col159[122] <= data_col159[121];
   data_col159[123] <= data_col159[122];
   data_col159[124] <= data_col159[123];
   data_col159[125] <= data_col159[124];
   data_col159[126] <= data_col159[125];
   data_col159[127] <= data_col159[126];
   data_col159[128] <= data_col159[127];
   data_col159[129] <= data_col159[128];
   data_col159[130] <= data_col159[129];
   data_col159[131] <= data_col159[130];
   data_col159[132] <= data_col159[131];
   data_col159[133] <= data_col159[132];
   data_col159[134] <= data_col159[133];
   data_col159[135] <= data_col159[134];
   data_col159[136] <= data_col159[135];
   data_col159[137] <= data_col159[136];
   data_col159[138] <= data_col159[137];
   data_col159[139] <= data_col159[138];
   data_col159[140] <= data_col159[139];
   data_col159[141] <= data_col159[140];
   data_col159[142] <= data_col159[141];
   data_col159[143] <= data_col159[142];
   data_col159[144] <= data_col159[143];
   data_col159[145] <= data_col159[144];
   data_col159[146] <= data_col159[145];
   data_col159[147] <= data_col159[146];
   data_col159[148] <= data_col159[147];
   data_col159[149] <= data_col159[148];
   data_col159[150] <= data_col159[149];
   data_col159[151] <= data_col159[150];
   data_col159[152] <= data_col159[151];
   data_col159[153] <= data_col159[152];
   data_col159[154] <= data_col159[153];
   data_col159[155] <= data_col159[154];
   data_col159[156] <= data_col159[155];
   data_col159[157] <= data_col159[156];
   data_col159[158] <= data_col159[157];
   data_col159[159] <= data_col159[158];

   data_col160[1] <= data[5];
   data_col160[2] <= data_col160[1];
   data_col160[3] <= data_col160[2];
   data_col160[4] <= data_col160[3];
   data_col160[5] <= data_col160[4];
   data_col160[6] <= data_col160[5];
   data_col160[7] <= data_col160[6];
   data_col160[8] <= data_col160[7];
   data_col160[9] <= data_col160[8];
   data_col160[10] <= data_col160[9];
   data_col160[11] <= data_col160[10];
   data_col160[12] <= data_col160[11];
   data_col160[13] <= data_col160[12];
   data_col160[14] <= data_col160[13];
   data_col160[15] <= data_col160[14];
   data_col160[16] <= data_col160[15];
   data_col160[17] <= data_col160[16];
   data_col160[18] <= data_col160[17];
   data_col160[19] <= data_col160[18];
   data_col160[20] <= data_col160[19];
   data_col160[21] <= data_col160[20];
   data_col160[22] <= data_col160[21];
   data_col160[23] <= data_col160[22];
   data_col160[24] <= data_col160[23];
   data_col160[25] <= data_col160[24];
   data_col160[26] <= data_col160[25];
   data_col160[27] <= data_col160[26];
   data_col160[28] <= data_col160[27];
   data_col160[29] <= data_col160[28];
   data_col160[30] <= data_col160[29];
   data_col160[31] <= data_col160[30];
   data_col160[32] <= data_col160[31];
   data_col160[33] <= data_col160[32];
   data_col160[34] <= data_col160[33];
   data_col160[35] <= data_col160[34];
   data_col160[36] <= data_col160[35];
   data_col160[37] <= data_col160[36];
   data_col160[38] <= data_col160[37];
   data_col160[39] <= data_col160[38];
   data_col160[40] <= data_col160[39];
   data_col160[41] <= data_col160[40];
   data_col160[42] <= data_col160[41];
   data_col160[43] <= data_col160[42];
   data_col160[44] <= data_col160[43];
   data_col160[45] <= data_col160[44];
   data_col160[46] <= data_col160[45];
   data_col160[47] <= data_col160[46];
   data_col160[48] <= data_col160[47];
   data_col160[49] <= data_col160[48];
   data_col160[50] <= data_col160[49];
   data_col160[51] <= data_col160[50];
   data_col160[52] <= data_col160[51];
   data_col160[53] <= data_col160[52];
   data_col160[54] <= data_col160[53];
   data_col160[55] <= data_col160[54];
   data_col160[56] <= data_col160[55];
   data_col160[57] <= data_col160[56];
   data_col160[58] <= data_col160[57];
   data_col160[59] <= data_col160[58];
   data_col160[60] <= data_col160[59];
   data_col160[61] <= data_col160[60];
   data_col160[62] <= data_col160[61];
   data_col160[63] <= data_col160[62];
   data_col160[64] <= data_col160[63];
   data_col160[65] <= data_col160[64];
   data_col160[66] <= data_col160[65];
   data_col160[67] <= data_col160[66];
   data_col160[68] <= data_col160[67];
   data_col160[69] <= data_col160[68];
   data_col160[70] <= data_col160[69];
   data_col160[71] <= data_col160[70];
   data_col160[72] <= data_col160[71];
   data_col160[73] <= data_col160[72];
   data_col160[74] <= data_col160[73];
   data_col160[75] <= data_col160[74];
   data_col160[76] <= data_col160[75];
   data_col160[77] <= data_col160[76];
   data_col160[78] <= data_col160[77];
   data_col160[79] <= data_col160[78];
   data_col160[80] <= data_col160[79];
   data_col160[81] <= data_col160[80];
   data_col160[82] <= data_col160[81];
   data_col160[83] <= data_col160[82];
   data_col160[84] <= data_col160[83];
   data_col160[85] <= data_col160[84];
   data_col160[86] <= data_col160[85];
   data_col160[87] <= data_col160[86];
   data_col160[88] <= data_col160[87];
   data_col160[89] <= data_col160[88];
   data_col160[90] <= data_col160[89];
   data_col160[91] <= data_col160[90];
   data_col160[92] <= data_col160[91];
   data_col160[93] <= data_col160[92];
   data_col160[94] <= data_col160[93];
   data_col160[95] <= data_col160[94];
   data_col160[96] <= data_col160[95];
   data_col160[97] <= data_col160[96];
   data_col160[98] <= data_col160[97];
   data_col160[99] <= data_col160[98];
   data_col160[100] <= data_col160[99];
   data_col160[101] <= data_col160[100];
   data_col160[102] <= data_col160[101];
   data_col160[103] <= data_col160[102];
   data_col160[104] <= data_col160[103];
   data_col160[105] <= data_col160[104];
   data_col160[106] <= data_col160[105];
   data_col160[107] <= data_col160[106];
   data_col160[108] <= data_col160[107];
   data_col160[109] <= data_col160[108];
   data_col160[110] <= data_col160[109];
   data_col160[111] <= data_col160[110];
   data_col160[112] <= data_col160[111];
   data_col160[113] <= data_col160[112];
   data_col160[114] <= data_col160[113];
   data_col160[115] <= data_col160[114];
   data_col160[116] <= data_col160[115];
   data_col160[117] <= data_col160[116];
   data_col160[118] <= data_col160[117];
   data_col160[119] <= data_col160[118];
   data_col160[120] <= data_col160[119];
   data_col160[121] <= data_col160[120];
   data_col160[122] <= data_col160[121];
   data_col160[123] <= data_col160[122];
   data_col160[124] <= data_col160[123];
   data_col160[125] <= data_col160[124];
   data_col160[126] <= data_col160[125];
   data_col160[127] <= data_col160[126];
   data_col160[128] <= data_col160[127];
   data_col160[129] <= data_col160[128];
   data_col160[130] <= data_col160[129];
   data_col160[131] <= data_col160[130];
   data_col160[132] <= data_col160[131];
   data_col160[133] <= data_col160[132];
   data_col160[134] <= data_col160[133];
   data_col160[135] <= data_col160[134];
   data_col160[136] <= data_col160[135];
   data_col160[137] <= data_col160[136];
   data_col160[138] <= data_col160[137];
   data_col160[139] <= data_col160[138];
   data_col160[140] <= data_col160[139];
   data_col160[141] <= data_col160[140];
   data_col160[142] <= data_col160[141];
   data_col160[143] <= data_col160[142];
   data_col160[144] <= data_col160[143];
   data_col160[145] <= data_col160[144];
   data_col160[146] <= data_col160[145];
   data_col160[147] <= data_col160[146];
   data_col160[148] <= data_col160[147];
   data_col160[149] <= data_col160[148];
   data_col160[150] <= data_col160[149];
   data_col160[151] <= data_col160[150];
   data_col160[152] <= data_col160[151];
   data_col160[153] <= data_col160[152];
   data_col160[154] <= data_col160[153];
   data_col160[155] <= data_col160[154];
   data_col160[156] <= data_col160[155];
   data_col160[157] <= data_col160[156];
   data_col160[158] <= data_col160[157];
   data_col160[159] <= data_col160[158];
   data_col160[160] <= data_col160[159];

   data_col161[1] <= data[4];
   data_col161[2] <= data_col161[1];
   data_col161[3] <= data_col161[2];
   data_col161[4] <= data_col161[3];
   data_col161[5] <= data_col161[4];
   data_col161[6] <= data_col161[5];
   data_col161[7] <= data_col161[6];
   data_col161[8] <= data_col161[7];
   data_col161[9] <= data_col161[8];
   data_col161[10] <= data_col161[9];
   data_col161[11] <= data_col161[10];
   data_col161[12] <= data_col161[11];
   data_col161[13] <= data_col161[12];
   data_col161[14] <= data_col161[13];
   data_col161[15] <= data_col161[14];
   data_col161[16] <= data_col161[15];
   data_col161[17] <= data_col161[16];
   data_col161[18] <= data_col161[17];
   data_col161[19] <= data_col161[18];
   data_col161[20] <= data_col161[19];
   data_col161[21] <= data_col161[20];
   data_col161[22] <= data_col161[21];
   data_col161[23] <= data_col161[22];
   data_col161[24] <= data_col161[23];
   data_col161[25] <= data_col161[24];
   data_col161[26] <= data_col161[25];
   data_col161[27] <= data_col161[26];
   data_col161[28] <= data_col161[27];
   data_col161[29] <= data_col161[28];
   data_col161[30] <= data_col161[29];
   data_col161[31] <= data_col161[30];
   data_col161[32] <= data_col161[31];
   data_col161[33] <= data_col161[32];
   data_col161[34] <= data_col161[33];
   data_col161[35] <= data_col161[34];
   data_col161[36] <= data_col161[35];
   data_col161[37] <= data_col161[36];
   data_col161[38] <= data_col161[37];
   data_col161[39] <= data_col161[38];
   data_col161[40] <= data_col161[39];
   data_col161[41] <= data_col161[40];
   data_col161[42] <= data_col161[41];
   data_col161[43] <= data_col161[42];
   data_col161[44] <= data_col161[43];
   data_col161[45] <= data_col161[44];
   data_col161[46] <= data_col161[45];
   data_col161[47] <= data_col161[46];
   data_col161[48] <= data_col161[47];
   data_col161[49] <= data_col161[48];
   data_col161[50] <= data_col161[49];
   data_col161[51] <= data_col161[50];
   data_col161[52] <= data_col161[51];
   data_col161[53] <= data_col161[52];
   data_col161[54] <= data_col161[53];
   data_col161[55] <= data_col161[54];
   data_col161[56] <= data_col161[55];
   data_col161[57] <= data_col161[56];
   data_col161[58] <= data_col161[57];
   data_col161[59] <= data_col161[58];
   data_col161[60] <= data_col161[59];
   data_col161[61] <= data_col161[60];
   data_col161[62] <= data_col161[61];
   data_col161[63] <= data_col161[62];
   data_col161[64] <= data_col161[63];
   data_col161[65] <= data_col161[64];
   data_col161[66] <= data_col161[65];
   data_col161[67] <= data_col161[66];
   data_col161[68] <= data_col161[67];
   data_col161[69] <= data_col161[68];
   data_col161[70] <= data_col161[69];
   data_col161[71] <= data_col161[70];
   data_col161[72] <= data_col161[71];
   data_col161[73] <= data_col161[72];
   data_col161[74] <= data_col161[73];
   data_col161[75] <= data_col161[74];
   data_col161[76] <= data_col161[75];
   data_col161[77] <= data_col161[76];
   data_col161[78] <= data_col161[77];
   data_col161[79] <= data_col161[78];
   data_col161[80] <= data_col161[79];
   data_col161[81] <= data_col161[80];
   data_col161[82] <= data_col161[81];
   data_col161[83] <= data_col161[82];
   data_col161[84] <= data_col161[83];
   data_col161[85] <= data_col161[84];
   data_col161[86] <= data_col161[85];
   data_col161[87] <= data_col161[86];
   data_col161[88] <= data_col161[87];
   data_col161[89] <= data_col161[88];
   data_col161[90] <= data_col161[89];
   data_col161[91] <= data_col161[90];
   data_col161[92] <= data_col161[91];
   data_col161[93] <= data_col161[92];
   data_col161[94] <= data_col161[93];
   data_col161[95] <= data_col161[94];
   data_col161[96] <= data_col161[95];
   data_col161[97] <= data_col161[96];
   data_col161[98] <= data_col161[97];
   data_col161[99] <= data_col161[98];
   data_col161[100] <= data_col161[99];
   data_col161[101] <= data_col161[100];
   data_col161[102] <= data_col161[101];
   data_col161[103] <= data_col161[102];
   data_col161[104] <= data_col161[103];
   data_col161[105] <= data_col161[104];
   data_col161[106] <= data_col161[105];
   data_col161[107] <= data_col161[106];
   data_col161[108] <= data_col161[107];
   data_col161[109] <= data_col161[108];
   data_col161[110] <= data_col161[109];
   data_col161[111] <= data_col161[110];
   data_col161[112] <= data_col161[111];
   data_col161[113] <= data_col161[112];
   data_col161[114] <= data_col161[113];
   data_col161[115] <= data_col161[114];
   data_col161[116] <= data_col161[115];
   data_col161[117] <= data_col161[116];
   data_col161[118] <= data_col161[117];
   data_col161[119] <= data_col161[118];
   data_col161[120] <= data_col161[119];
   data_col161[121] <= data_col161[120];
   data_col161[122] <= data_col161[121];
   data_col161[123] <= data_col161[122];
   data_col161[124] <= data_col161[123];
   data_col161[125] <= data_col161[124];
   data_col161[126] <= data_col161[125];
   data_col161[127] <= data_col161[126];
   data_col161[128] <= data_col161[127];
   data_col161[129] <= data_col161[128];
   data_col161[130] <= data_col161[129];
   data_col161[131] <= data_col161[130];
   data_col161[132] <= data_col161[131];
   data_col161[133] <= data_col161[132];
   data_col161[134] <= data_col161[133];
   data_col161[135] <= data_col161[134];
   data_col161[136] <= data_col161[135];
   data_col161[137] <= data_col161[136];
   data_col161[138] <= data_col161[137];
   data_col161[139] <= data_col161[138];
   data_col161[140] <= data_col161[139];
   data_col161[141] <= data_col161[140];
   data_col161[142] <= data_col161[141];
   data_col161[143] <= data_col161[142];
   data_col161[144] <= data_col161[143];
   data_col161[145] <= data_col161[144];
   data_col161[146] <= data_col161[145];
   data_col161[147] <= data_col161[146];
   data_col161[148] <= data_col161[147];
   data_col161[149] <= data_col161[148];
   data_col161[150] <= data_col161[149];
   data_col161[151] <= data_col161[150];
   data_col161[152] <= data_col161[151];
   data_col161[153] <= data_col161[152];
   data_col161[154] <= data_col161[153];
   data_col161[155] <= data_col161[154];
   data_col161[156] <= data_col161[155];
   data_col161[157] <= data_col161[156];
   data_col161[158] <= data_col161[157];
   data_col161[159] <= data_col161[158];
   data_col161[160] <= data_col161[159];
   data_col161[161] <= data_col161[160];

   data_col162[1] <= data[3];
   data_col162[2] <= data_col162[1];
   data_col162[3] <= data_col162[2];
   data_col162[4] <= data_col162[3];
   data_col162[5] <= data_col162[4];
   data_col162[6] <= data_col162[5];
   data_col162[7] <= data_col162[6];
   data_col162[8] <= data_col162[7];
   data_col162[9] <= data_col162[8];
   data_col162[10] <= data_col162[9];
   data_col162[11] <= data_col162[10];
   data_col162[12] <= data_col162[11];
   data_col162[13] <= data_col162[12];
   data_col162[14] <= data_col162[13];
   data_col162[15] <= data_col162[14];
   data_col162[16] <= data_col162[15];
   data_col162[17] <= data_col162[16];
   data_col162[18] <= data_col162[17];
   data_col162[19] <= data_col162[18];
   data_col162[20] <= data_col162[19];
   data_col162[21] <= data_col162[20];
   data_col162[22] <= data_col162[21];
   data_col162[23] <= data_col162[22];
   data_col162[24] <= data_col162[23];
   data_col162[25] <= data_col162[24];
   data_col162[26] <= data_col162[25];
   data_col162[27] <= data_col162[26];
   data_col162[28] <= data_col162[27];
   data_col162[29] <= data_col162[28];
   data_col162[30] <= data_col162[29];
   data_col162[31] <= data_col162[30];
   data_col162[32] <= data_col162[31];
   data_col162[33] <= data_col162[32];
   data_col162[34] <= data_col162[33];
   data_col162[35] <= data_col162[34];
   data_col162[36] <= data_col162[35];
   data_col162[37] <= data_col162[36];
   data_col162[38] <= data_col162[37];
   data_col162[39] <= data_col162[38];
   data_col162[40] <= data_col162[39];
   data_col162[41] <= data_col162[40];
   data_col162[42] <= data_col162[41];
   data_col162[43] <= data_col162[42];
   data_col162[44] <= data_col162[43];
   data_col162[45] <= data_col162[44];
   data_col162[46] <= data_col162[45];
   data_col162[47] <= data_col162[46];
   data_col162[48] <= data_col162[47];
   data_col162[49] <= data_col162[48];
   data_col162[50] <= data_col162[49];
   data_col162[51] <= data_col162[50];
   data_col162[52] <= data_col162[51];
   data_col162[53] <= data_col162[52];
   data_col162[54] <= data_col162[53];
   data_col162[55] <= data_col162[54];
   data_col162[56] <= data_col162[55];
   data_col162[57] <= data_col162[56];
   data_col162[58] <= data_col162[57];
   data_col162[59] <= data_col162[58];
   data_col162[60] <= data_col162[59];
   data_col162[61] <= data_col162[60];
   data_col162[62] <= data_col162[61];
   data_col162[63] <= data_col162[62];
   data_col162[64] <= data_col162[63];
   data_col162[65] <= data_col162[64];
   data_col162[66] <= data_col162[65];
   data_col162[67] <= data_col162[66];
   data_col162[68] <= data_col162[67];
   data_col162[69] <= data_col162[68];
   data_col162[70] <= data_col162[69];
   data_col162[71] <= data_col162[70];
   data_col162[72] <= data_col162[71];
   data_col162[73] <= data_col162[72];
   data_col162[74] <= data_col162[73];
   data_col162[75] <= data_col162[74];
   data_col162[76] <= data_col162[75];
   data_col162[77] <= data_col162[76];
   data_col162[78] <= data_col162[77];
   data_col162[79] <= data_col162[78];
   data_col162[80] <= data_col162[79];
   data_col162[81] <= data_col162[80];
   data_col162[82] <= data_col162[81];
   data_col162[83] <= data_col162[82];
   data_col162[84] <= data_col162[83];
   data_col162[85] <= data_col162[84];
   data_col162[86] <= data_col162[85];
   data_col162[87] <= data_col162[86];
   data_col162[88] <= data_col162[87];
   data_col162[89] <= data_col162[88];
   data_col162[90] <= data_col162[89];
   data_col162[91] <= data_col162[90];
   data_col162[92] <= data_col162[91];
   data_col162[93] <= data_col162[92];
   data_col162[94] <= data_col162[93];
   data_col162[95] <= data_col162[94];
   data_col162[96] <= data_col162[95];
   data_col162[97] <= data_col162[96];
   data_col162[98] <= data_col162[97];
   data_col162[99] <= data_col162[98];
   data_col162[100] <= data_col162[99];
   data_col162[101] <= data_col162[100];
   data_col162[102] <= data_col162[101];
   data_col162[103] <= data_col162[102];
   data_col162[104] <= data_col162[103];
   data_col162[105] <= data_col162[104];
   data_col162[106] <= data_col162[105];
   data_col162[107] <= data_col162[106];
   data_col162[108] <= data_col162[107];
   data_col162[109] <= data_col162[108];
   data_col162[110] <= data_col162[109];
   data_col162[111] <= data_col162[110];
   data_col162[112] <= data_col162[111];
   data_col162[113] <= data_col162[112];
   data_col162[114] <= data_col162[113];
   data_col162[115] <= data_col162[114];
   data_col162[116] <= data_col162[115];
   data_col162[117] <= data_col162[116];
   data_col162[118] <= data_col162[117];
   data_col162[119] <= data_col162[118];
   data_col162[120] <= data_col162[119];
   data_col162[121] <= data_col162[120];
   data_col162[122] <= data_col162[121];
   data_col162[123] <= data_col162[122];
   data_col162[124] <= data_col162[123];
   data_col162[125] <= data_col162[124];
   data_col162[126] <= data_col162[125];
   data_col162[127] <= data_col162[126];
   data_col162[128] <= data_col162[127];
   data_col162[129] <= data_col162[128];
   data_col162[130] <= data_col162[129];
   data_col162[131] <= data_col162[130];
   data_col162[132] <= data_col162[131];
   data_col162[133] <= data_col162[132];
   data_col162[134] <= data_col162[133];
   data_col162[135] <= data_col162[134];
   data_col162[136] <= data_col162[135];
   data_col162[137] <= data_col162[136];
   data_col162[138] <= data_col162[137];
   data_col162[139] <= data_col162[138];
   data_col162[140] <= data_col162[139];
   data_col162[141] <= data_col162[140];
   data_col162[142] <= data_col162[141];
   data_col162[143] <= data_col162[142];
   data_col162[144] <= data_col162[143];
   data_col162[145] <= data_col162[144];
   data_col162[146] <= data_col162[145];
   data_col162[147] <= data_col162[146];
   data_col162[148] <= data_col162[147];
   data_col162[149] <= data_col162[148];
   data_col162[150] <= data_col162[149];
   data_col162[151] <= data_col162[150];
   data_col162[152] <= data_col162[151];
   data_col162[153] <= data_col162[152];
   data_col162[154] <= data_col162[153];
   data_col162[155] <= data_col162[154];
   data_col162[156] <= data_col162[155];
   data_col162[157] <= data_col162[156];
   data_col162[158] <= data_col162[157];
   data_col162[159] <= data_col162[158];
   data_col162[160] <= data_col162[159];
   data_col162[161] <= data_col162[160];
   data_col162[162] <= data_col162[161];

   data_col163[1] <= data[2];
   data_col163[2] <= data_col163[1];
   data_col163[3] <= data_col163[2];
   data_col163[4] <= data_col163[3];
   data_col163[5] <= data_col163[4];
   data_col163[6] <= data_col163[5];
   data_col163[7] <= data_col163[6];
   data_col163[8] <= data_col163[7];
   data_col163[9] <= data_col163[8];
   data_col163[10] <= data_col163[9];
   data_col163[11] <= data_col163[10];
   data_col163[12] <= data_col163[11];
   data_col163[13] <= data_col163[12];
   data_col163[14] <= data_col163[13];
   data_col163[15] <= data_col163[14];
   data_col163[16] <= data_col163[15];
   data_col163[17] <= data_col163[16];
   data_col163[18] <= data_col163[17];
   data_col163[19] <= data_col163[18];
   data_col163[20] <= data_col163[19];
   data_col163[21] <= data_col163[20];
   data_col163[22] <= data_col163[21];
   data_col163[23] <= data_col163[22];
   data_col163[24] <= data_col163[23];
   data_col163[25] <= data_col163[24];
   data_col163[26] <= data_col163[25];
   data_col163[27] <= data_col163[26];
   data_col163[28] <= data_col163[27];
   data_col163[29] <= data_col163[28];
   data_col163[30] <= data_col163[29];
   data_col163[31] <= data_col163[30];
   data_col163[32] <= data_col163[31];
   data_col163[33] <= data_col163[32];
   data_col163[34] <= data_col163[33];
   data_col163[35] <= data_col163[34];
   data_col163[36] <= data_col163[35];
   data_col163[37] <= data_col163[36];
   data_col163[38] <= data_col163[37];
   data_col163[39] <= data_col163[38];
   data_col163[40] <= data_col163[39];
   data_col163[41] <= data_col163[40];
   data_col163[42] <= data_col163[41];
   data_col163[43] <= data_col163[42];
   data_col163[44] <= data_col163[43];
   data_col163[45] <= data_col163[44];
   data_col163[46] <= data_col163[45];
   data_col163[47] <= data_col163[46];
   data_col163[48] <= data_col163[47];
   data_col163[49] <= data_col163[48];
   data_col163[50] <= data_col163[49];
   data_col163[51] <= data_col163[50];
   data_col163[52] <= data_col163[51];
   data_col163[53] <= data_col163[52];
   data_col163[54] <= data_col163[53];
   data_col163[55] <= data_col163[54];
   data_col163[56] <= data_col163[55];
   data_col163[57] <= data_col163[56];
   data_col163[58] <= data_col163[57];
   data_col163[59] <= data_col163[58];
   data_col163[60] <= data_col163[59];
   data_col163[61] <= data_col163[60];
   data_col163[62] <= data_col163[61];
   data_col163[63] <= data_col163[62];
   data_col163[64] <= data_col163[63];
   data_col163[65] <= data_col163[64];
   data_col163[66] <= data_col163[65];
   data_col163[67] <= data_col163[66];
   data_col163[68] <= data_col163[67];
   data_col163[69] <= data_col163[68];
   data_col163[70] <= data_col163[69];
   data_col163[71] <= data_col163[70];
   data_col163[72] <= data_col163[71];
   data_col163[73] <= data_col163[72];
   data_col163[74] <= data_col163[73];
   data_col163[75] <= data_col163[74];
   data_col163[76] <= data_col163[75];
   data_col163[77] <= data_col163[76];
   data_col163[78] <= data_col163[77];
   data_col163[79] <= data_col163[78];
   data_col163[80] <= data_col163[79];
   data_col163[81] <= data_col163[80];
   data_col163[82] <= data_col163[81];
   data_col163[83] <= data_col163[82];
   data_col163[84] <= data_col163[83];
   data_col163[85] <= data_col163[84];
   data_col163[86] <= data_col163[85];
   data_col163[87] <= data_col163[86];
   data_col163[88] <= data_col163[87];
   data_col163[89] <= data_col163[88];
   data_col163[90] <= data_col163[89];
   data_col163[91] <= data_col163[90];
   data_col163[92] <= data_col163[91];
   data_col163[93] <= data_col163[92];
   data_col163[94] <= data_col163[93];
   data_col163[95] <= data_col163[94];
   data_col163[96] <= data_col163[95];
   data_col163[97] <= data_col163[96];
   data_col163[98] <= data_col163[97];
   data_col163[99] <= data_col163[98];
   data_col163[100] <= data_col163[99];
   data_col163[101] <= data_col163[100];
   data_col163[102] <= data_col163[101];
   data_col163[103] <= data_col163[102];
   data_col163[104] <= data_col163[103];
   data_col163[105] <= data_col163[104];
   data_col163[106] <= data_col163[105];
   data_col163[107] <= data_col163[106];
   data_col163[108] <= data_col163[107];
   data_col163[109] <= data_col163[108];
   data_col163[110] <= data_col163[109];
   data_col163[111] <= data_col163[110];
   data_col163[112] <= data_col163[111];
   data_col163[113] <= data_col163[112];
   data_col163[114] <= data_col163[113];
   data_col163[115] <= data_col163[114];
   data_col163[116] <= data_col163[115];
   data_col163[117] <= data_col163[116];
   data_col163[118] <= data_col163[117];
   data_col163[119] <= data_col163[118];
   data_col163[120] <= data_col163[119];
   data_col163[121] <= data_col163[120];
   data_col163[122] <= data_col163[121];
   data_col163[123] <= data_col163[122];
   data_col163[124] <= data_col163[123];
   data_col163[125] <= data_col163[124];
   data_col163[126] <= data_col163[125];
   data_col163[127] <= data_col163[126];
   data_col163[128] <= data_col163[127];
   data_col163[129] <= data_col163[128];
   data_col163[130] <= data_col163[129];
   data_col163[131] <= data_col163[130];
   data_col163[132] <= data_col163[131];
   data_col163[133] <= data_col163[132];
   data_col163[134] <= data_col163[133];
   data_col163[135] <= data_col163[134];
   data_col163[136] <= data_col163[135];
   data_col163[137] <= data_col163[136];
   data_col163[138] <= data_col163[137];
   data_col163[139] <= data_col163[138];
   data_col163[140] <= data_col163[139];
   data_col163[141] <= data_col163[140];
   data_col163[142] <= data_col163[141];
   data_col163[143] <= data_col163[142];
   data_col163[144] <= data_col163[143];
   data_col163[145] <= data_col163[144];
   data_col163[146] <= data_col163[145];
   data_col163[147] <= data_col163[146];
   data_col163[148] <= data_col163[147];
   data_col163[149] <= data_col163[148];
   data_col163[150] <= data_col163[149];
   data_col163[151] <= data_col163[150];
   data_col163[152] <= data_col163[151];
   data_col163[153] <= data_col163[152];
   data_col163[154] <= data_col163[153];
   data_col163[155] <= data_col163[154];
   data_col163[156] <= data_col163[155];
   data_col163[157] <= data_col163[156];
   data_col163[158] <= data_col163[157];
   data_col163[159] <= data_col163[158];
   data_col163[160] <= data_col163[159];
   data_col163[161] <= data_col163[160];
   data_col163[162] <= data_col163[161];
   data_col163[163] <= data_col163[162];

   data_col164[1] <= data[1];
   data_col164[2] <= data_col164[1];
   data_col164[3] <= data_col164[2];
   data_col164[4] <= data_col164[3];
   data_col164[5] <= data_col164[4];
   data_col164[6] <= data_col164[5];
   data_col164[7] <= data_col164[6];
   data_col164[8] <= data_col164[7];
   data_col164[9] <= data_col164[8];
   data_col164[10] <= data_col164[9];
   data_col164[11] <= data_col164[10];
   data_col164[12] <= data_col164[11];
   data_col164[13] <= data_col164[12];
   data_col164[14] <= data_col164[13];
   data_col164[15] <= data_col164[14];
   data_col164[16] <= data_col164[15];
   data_col164[17] <= data_col164[16];
   data_col164[18] <= data_col164[17];
   data_col164[19] <= data_col164[18];
   data_col164[20] <= data_col164[19];
   data_col164[21] <= data_col164[20];
   data_col164[22] <= data_col164[21];
   data_col164[23] <= data_col164[22];
   data_col164[24] <= data_col164[23];
   data_col164[25] <= data_col164[24];
   data_col164[26] <= data_col164[25];
   data_col164[27] <= data_col164[26];
   data_col164[28] <= data_col164[27];
   data_col164[29] <= data_col164[28];
   data_col164[30] <= data_col164[29];
   data_col164[31] <= data_col164[30];
   data_col164[32] <= data_col164[31];
   data_col164[33] <= data_col164[32];
   data_col164[34] <= data_col164[33];
   data_col164[35] <= data_col164[34];
   data_col164[36] <= data_col164[35];
   data_col164[37] <= data_col164[36];
   data_col164[38] <= data_col164[37];
   data_col164[39] <= data_col164[38];
   data_col164[40] <= data_col164[39];
   data_col164[41] <= data_col164[40];
   data_col164[42] <= data_col164[41];
   data_col164[43] <= data_col164[42];
   data_col164[44] <= data_col164[43];
   data_col164[45] <= data_col164[44];
   data_col164[46] <= data_col164[45];
   data_col164[47] <= data_col164[46];
   data_col164[48] <= data_col164[47];
   data_col164[49] <= data_col164[48];
   data_col164[50] <= data_col164[49];
   data_col164[51] <= data_col164[50];
   data_col164[52] <= data_col164[51];
   data_col164[53] <= data_col164[52];
   data_col164[54] <= data_col164[53];
   data_col164[55] <= data_col164[54];
   data_col164[56] <= data_col164[55];
   data_col164[57] <= data_col164[56];
   data_col164[58] <= data_col164[57];
   data_col164[59] <= data_col164[58];
   data_col164[60] <= data_col164[59];
   data_col164[61] <= data_col164[60];
   data_col164[62] <= data_col164[61];
   data_col164[63] <= data_col164[62];
   data_col164[64] <= data_col164[63];
   data_col164[65] <= data_col164[64];
   data_col164[66] <= data_col164[65];
   data_col164[67] <= data_col164[66];
   data_col164[68] <= data_col164[67];
   data_col164[69] <= data_col164[68];
   data_col164[70] <= data_col164[69];
   data_col164[71] <= data_col164[70];
   data_col164[72] <= data_col164[71];
   data_col164[73] <= data_col164[72];
   data_col164[74] <= data_col164[73];
   data_col164[75] <= data_col164[74];
   data_col164[76] <= data_col164[75];
   data_col164[77] <= data_col164[76];
   data_col164[78] <= data_col164[77];
   data_col164[79] <= data_col164[78];
   data_col164[80] <= data_col164[79];
   data_col164[81] <= data_col164[80];
   data_col164[82] <= data_col164[81];
   data_col164[83] <= data_col164[82];
   data_col164[84] <= data_col164[83];
   data_col164[85] <= data_col164[84];
   data_col164[86] <= data_col164[85];
   data_col164[87] <= data_col164[86];
   data_col164[88] <= data_col164[87];
   data_col164[89] <= data_col164[88];
   data_col164[90] <= data_col164[89];
   data_col164[91] <= data_col164[90];
   data_col164[92] <= data_col164[91];
   data_col164[93] <= data_col164[92];
   data_col164[94] <= data_col164[93];
   data_col164[95] <= data_col164[94];
   data_col164[96] <= data_col164[95];
   data_col164[97] <= data_col164[96];
   data_col164[98] <= data_col164[97];
   data_col164[99] <= data_col164[98];
   data_col164[100] <= data_col164[99];
   data_col164[101] <= data_col164[100];
   data_col164[102] <= data_col164[101];
   data_col164[103] <= data_col164[102];
   data_col164[104] <= data_col164[103];
   data_col164[105] <= data_col164[104];
   data_col164[106] <= data_col164[105];
   data_col164[107] <= data_col164[106];
   data_col164[108] <= data_col164[107];
   data_col164[109] <= data_col164[108];
   data_col164[110] <= data_col164[109];
   data_col164[111] <= data_col164[110];
   data_col164[112] <= data_col164[111];
   data_col164[113] <= data_col164[112];
   data_col164[114] <= data_col164[113];
   data_col164[115] <= data_col164[114];
   data_col164[116] <= data_col164[115];
   data_col164[117] <= data_col164[116];
   data_col164[118] <= data_col164[117];
   data_col164[119] <= data_col164[118];
   data_col164[120] <= data_col164[119];
   data_col164[121] <= data_col164[120];
   data_col164[122] <= data_col164[121];
   data_col164[123] <= data_col164[122];
   data_col164[124] <= data_col164[123];
   data_col164[125] <= data_col164[124];
   data_col164[126] <= data_col164[125];
   data_col164[127] <= data_col164[126];
   data_col164[128] <= data_col164[127];
   data_col164[129] <= data_col164[128];
   data_col164[130] <= data_col164[129];
   data_col164[131] <= data_col164[130];
   data_col164[132] <= data_col164[131];
   data_col164[133] <= data_col164[132];
   data_col164[134] <= data_col164[133];
   data_col164[135] <= data_col164[134];
   data_col164[136] <= data_col164[135];
   data_col164[137] <= data_col164[136];
   data_col164[138] <= data_col164[137];
   data_col164[139] <= data_col164[138];
   data_col164[140] <= data_col164[139];
   data_col164[141] <= data_col164[140];
   data_col164[142] <= data_col164[141];
   data_col164[143] <= data_col164[142];
   data_col164[144] <= data_col164[143];
   data_col164[145] <= data_col164[144];
   data_col164[146] <= data_col164[145];
   data_col164[147] <= data_col164[146];
   data_col164[148] <= data_col164[147];
   data_col164[149] <= data_col164[148];
   data_col164[150] <= data_col164[149];
   data_col164[151] <= data_col164[150];
   data_col164[152] <= data_col164[151];
   data_col164[153] <= data_col164[152];
   data_col164[154] <= data_col164[153];
   data_col164[155] <= data_col164[154];
   data_col164[156] <= data_col164[155];
   data_col164[157] <= data_col164[156];
   data_col164[158] <= data_col164[157];
   data_col164[159] <= data_col164[158];
   data_col164[160] <= data_col164[159];
   data_col164[161] <= data_col164[160];
   data_col164[162] <= data_col164[161];
   data_col164[163] <= data_col164[162];
   data_col164[164] <= data_col164[163];

   data_col165[1] <= data[0];
   data_col165[2] <= data_col165[1];
   data_col165[3] <= data_col165[2];
   data_col165[4] <= data_col165[3];
   data_col165[5] <= data_col165[4];
   data_col165[6] <= data_col165[5];
   data_col165[7] <= data_col165[6];
   data_col165[8] <= data_col165[7];
   data_col165[9] <= data_col165[8];
   data_col165[10] <= data_col165[9];
   data_col165[11] <= data_col165[10];
   data_col165[12] <= data_col165[11];
   data_col165[13] <= data_col165[12];
   data_col165[14] <= data_col165[13];
   data_col165[15] <= data_col165[14];
   data_col165[16] <= data_col165[15];
   data_col165[17] <= data_col165[16];
   data_col165[18] <= data_col165[17];
   data_col165[19] <= data_col165[18];
   data_col165[20] <= data_col165[19];
   data_col165[21] <= data_col165[20];
   data_col165[22] <= data_col165[21];
   data_col165[23] <= data_col165[22];
   data_col165[24] <= data_col165[23];
   data_col165[25] <= data_col165[24];
   data_col165[26] <= data_col165[25];
   data_col165[27] <= data_col165[26];
   data_col165[28] <= data_col165[27];
   data_col165[29] <= data_col165[28];
   data_col165[30] <= data_col165[29];
   data_col165[31] <= data_col165[30];
   data_col165[32] <= data_col165[31];
   data_col165[33] <= data_col165[32];
   data_col165[34] <= data_col165[33];
   data_col165[35] <= data_col165[34];
   data_col165[36] <= data_col165[35];
   data_col165[37] <= data_col165[36];
   data_col165[38] <= data_col165[37];
   data_col165[39] <= data_col165[38];
   data_col165[40] <= data_col165[39];
   data_col165[41] <= data_col165[40];
   data_col165[42] <= data_col165[41];
   data_col165[43] <= data_col165[42];
   data_col165[44] <= data_col165[43];
   data_col165[45] <= data_col165[44];
   data_col165[46] <= data_col165[45];
   data_col165[47] <= data_col165[46];
   data_col165[48] <= data_col165[47];
   data_col165[49] <= data_col165[48];
   data_col165[50] <= data_col165[49];
   data_col165[51] <= data_col165[50];
   data_col165[52] <= data_col165[51];
   data_col165[53] <= data_col165[52];
   data_col165[54] <= data_col165[53];
   data_col165[55] <= data_col165[54];
   data_col165[56] <= data_col165[55];
   data_col165[57] <= data_col165[56];
   data_col165[58] <= data_col165[57];
   data_col165[59] <= data_col165[58];
   data_col165[60] <= data_col165[59];
   data_col165[61] <= data_col165[60];
   data_col165[62] <= data_col165[61];
   data_col165[63] <= data_col165[62];
   data_col165[64] <= data_col165[63];
   data_col165[65] <= data_col165[64];
   data_col165[66] <= data_col165[65];
   data_col165[67] <= data_col165[66];
   data_col165[68] <= data_col165[67];
   data_col165[69] <= data_col165[68];
   data_col165[70] <= data_col165[69];
   data_col165[71] <= data_col165[70];
   data_col165[72] <= data_col165[71];
   data_col165[73] <= data_col165[72];
   data_col165[74] <= data_col165[73];
   data_col165[75] <= data_col165[74];
   data_col165[76] <= data_col165[75];
   data_col165[77] <= data_col165[76];
   data_col165[78] <= data_col165[77];
   data_col165[79] <= data_col165[78];
   data_col165[80] <= data_col165[79];
   data_col165[81] <= data_col165[80];
   data_col165[82] <= data_col165[81];
   data_col165[83] <= data_col165[82];
   data_col165[84] <= data_col165[83];
   data_col165[85] <= data_col165[84];
   data_col165[86] <= data_col165[85];
   data_col165[87] <= data_col165[86];
   data_col165[88] <= data_col165[87];
   data_col165[89] <= data_col165[88];
   data_col165[90] <= data_col165[89];
   data_col165[91] <= data_col165[90];
   data_col165[92] <= data_col165[91];
   data_col165[93] <= data_col165[92];
   data_col165[94] <= data_col165[93];
   data_col165[95] <= data_col165[94];
   data_col165[96] <= data_col165[95];
   data_col165[97] <= data_col165[96];
   data_col165[98] <= data_col165[97];
   data_col165[99] <= data_col165[98];
   data_col165[100] <= data_col165[99];
   data_col165[101] <= data_col165[100];
   data_col165[102] <= data_col165[101];
   data_col165[103] <= data_col165[102];
   data_col165[104] <= data_col165[103];
   data_col165[105] <= data_col165[104];
   data_col165[106] <= data_col165[105];
   data_col165[107] <= data_col165[106];
   data_col165[108] <= data_col165[107];
   data_col165[109] <= data_col165[108];
   data_col165[110] <= data_col165[109];
   data_col165[111] <= data_col165[110];
   data_col165[112] <= data_col165[111];
   data_col165[113] <= data_col165[112];
   data_col165[114] <= data_col165[113];
   data_col165[115] <= data_col165[114];
   data_col165[116] <= data_col165[115];
   data_col165[117] <= data_col165[116];
   data_col165[118] <= data_col165[117];
   data_col165[119] <= data_col165[118];
   data_col165[120] <= data_col165[119];
   data_col165[121] <= data_col165[120];
   data_col165[122] <= data_col165[121];
   data_col165[123] <= data_col165[122];
   data_col165[124] <= data_col165[123];
   data_col165[125] <= data_col165[124];
   data_col165[126] <= data_col165[125];
   data_col165[127] <= data_col165[126];
   data_col165[128] <= data_col165[127];
   data_col165[129] <= data_col165[128];
   data_col165[130] <= data_col165[129];
   data_col165[131] <= data_col165[130];
   data_col165[132] <= data_col165[131];
   data_col165[133] <= data_col165[132];
   data_col165[134] <= data_col165[133];
   data_col165[135] <= data_col165[134];
   data_col165[136] <= data_col165[135];
   data_col165[137] <= data_col165[136];
   data_col165[138] <= data_col165[137];
   data_col165[139] <= data_col165[138];
   data_col165[140] <= data_col165[139];
   data_col165[141] <= data_col165[140];
   data_col165[142] <= data_col165[141];
   data_col165[143] <= data_col165[142];
   data_col165[144] <= data_col165[143];
   data_col165[145] <= data_col165[144];
   data_col165[146] <= data_col165[145];
   data_col165[147] <= data_col165[146];
   data_col165[148] <= data_col165[147];
   data_col165[149] <= data_col165[148];
   data_col165[150] <= data_col165[149];
   data_col165[151] <= data_col165[150];
   data_col165[152] <= data_col165[151];
   data_col165[153] <= data_col165[152];
   data_col165[154] <= data_col165[153];
   data_col165[155] <= data_col165[154];
   data_col165[156] <= data_col165[155];
   data_col165[157] <= data_col165[156];
   data_col165[158] <= data_col165[157];
   data_col165[159] <= data_col165[158];
   data_col165[160] <= data_col165[159];
   data_col165[161] <= data_col165[160];
   data_col165[162] <= data_col165[161];
   data_col165[163] <= data_col165[162];
   data_col165[164] <= data_col165[163];
   data_col165[165] <= data_col165[164];
 end

 wire [DAT_W-1:0] data_in;
 assign data_in = {data_col0, data_col1[1], data_col2[2], data_col3[3], data_col4[4], data_col5[5], data_col6[6], data_col7[7], data_col8[8], data_col9[9], data_col10[10], data_col11[11], data_col12[12], data_col13[13], data_col14[14], data_col15[15], data_col16[16], data_col17[17], data_col18[18], data_col19[19], data_col20[20], data_col21[21], data_col22[22], data_col23[23], data_col24[24], data_col25[25], data_col26[26], data_col27[27], data_col28[28], data_col29[29], data_col30[30], data_col31[31], data_col32[32], data_col33[33], data_col34[34], data_col35[35], data_col36[36], data_col37[37], data_col38[38], data_col39[39], data_col40[40], data_col41[41], data_col42[42], data_col43[43], data_col44[44], data_col45[45], data_col46[46], data_col47[47], data_col48[48], data_col49[49], data_col50[50], data_col51[51], data_col52[52], data_col53[53], data_col54[54], data_col55[55], data_col56[56], data_col57[57], data_col58[58], data_col59[59], data_col60[60], data_col61[61], data_col62[62], data_col63[63], data_col64[64], data_col65[65], data_col66[66], data_col67[67], data_col68[68], data_col69[69], data_col70[70], data_col71[71], data_col72[72], data_col73[73], data_col74[74], data_col75[75], data_col76[76], data_col77[77], data_col78[78], data_col79[79], data_col80[80], data_col81[81], data_col82[82], data_col83[83], data_col84[84], data_col85[85], data_col86[86], data_col87[87], data_col88[88], data_col89[89], data_col90[90], data_col91[91], data_col92[92], data_col93[93], data_col94[94], data_col95[95], data_col96[96], data_col97[97], data_col98[98], data_col99[99], data_col100[100], data_col101[101], data_col102[102], data_col103[103], data_col104[104], data_col105[105], data_col106[106], data_col107[107], data_col108[108], data_col109[109], data_col110[110], data_col111[111], data_col112[112], data_col113[113], data_col114[114], data_col115[115], data_col116[116], data_col117[117], data_col118[118], data_col119[119], data_col120[120], data_col121[121], data_col122[122], data_col123[123], data_col124[124], data_col125[125], data_col126[126], data_col127[127], data_col128[128], data_col129[129], data_col130[130], data_col131[131], data_col132[132], data_col133[133], data_col134[134], data_col135[135], data_col136[136], data_col137[137], data_col138[138], data_col139[139], data_col140[140], data_col141[141], data_col142[142], data_col143[143], data_col144[144], data_col145[145], data_col146[146], data_col147[147], data_col148[148], data_col149[149], data_col150[150], data_col151[151], data_col152[152], data_col153[153], data_col154[154], data_col155[155], data_col156[156], data_col157[157], data_col158[158], data_col159[159], data_col160[160], data_col161[161], data_col162[162], data_col163[163], data_col164[164], data_col165[165]};

  /////////////////////////////////////
  // row 0
  // row 0, col 0

     wire start_in_0_0;
     wire start_out_0_0;

     wire swap_in_0_0;
     wire swap_out_0_0;

     wire [1:0] op_in_0_0;
     wire [1:0] op_out_0_0;

     wire r_0_0;

     wire data_in_0_0;
     wire data_out_0_0;

     wire pivot_in_0_0;
     wire pivot_out_0_0;

     assign data_in_0_0 = data_in[DAT_W-1];
     assign op_in_0_0 = 2'b00;
     assign pivot_in_0_0 = 0;

     assign start_in_0_0 = start;
     assign swap_in_0_0 = swap;

     processor_AB AB_0_0 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_0),
       .start_in   (start_in_0_0),
       .swap_in    (swap_in_0_0),
       .op_in      (op_in_0_0),
       .pivot_in   (pivot_in_0_0),
       .start_out  (start_out_0_0),
       .swap_out   (swap_out_0_0),
       .data_out   (data_out_0_0),
       .op_out     (op_out_0_0),
       .pivot_out  (pivot_out_0_0),
       .r          (r_0_0)
     );

  // row 0, col 1

     reg start_in_0_1;
     wire start_out_0_1;

     reg swap_in_0_1;
     wire swap_out_0_1;

     reg [1:0] op_in_0_1;
     wire [1:0] op_out_0_1;

     wire r_0_1;

     wire data_in_0_1;
     wire data_out_0_1;

     reg pivot_in_0_1;
     wire pivot_out_0_1;

     assign data_in_0_1 = data_in[DAT_W-2];

     always @(posedge clk) begin
        op_in_0_1 <= op_out_0_0;
        pivot_in_0_1 <= pivot_out_0_0;
        start_in_0_1 <= start_out_0_0;
        swap_in_0_1 <= swap_out_0_0;
     end
  
     processor_AB AB_0_1 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_1),
       .start_in   (start_in_0_1),
       .swap_in    (swap_in_0_1),
       .op_in      (op_in_0_1),
       .pivot_in   (pivot_in_0_1),
       .start_out  (start_out_0_1),
       .swap_out   (swap_out_0_1),
       .data_out   (data_out_0_1),
       .op_out     (op_out_0_1),
       .pivot_out  (pivot_out_0_1),
       .r          (r_0_1)
     );

  // row 0, col 2

     reg start_in_0_2;
     wire start_out_0_2;

     reg swap_in_0_2;
     wire swap_out_0_2;

     reg [1:0] op_in_0_2;
     wire [1:0] op_out_0_2;

     wire r_0_2;

     wire data_in_0_2;
     wire data_out_0_2;

     reg pivot_in_0_2;
     wire pivot_out_0_2;

     assign data_in_0_2 = data_in[DAT_W-3];

     always @(posedge clk) begin
        op_in_0_2 <= op_out_0_1;
        pivot_in_0_2 <= pivot_out_0_1;
        start_in_0_2 <= start_out_0_1;
        swap_in_0_2 <= swap_out_0_1;
     end
  
     processor_AB AB_0_2 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_2),
       .start_in   (start_in_0_2),
       .swap_in    (swap_in_0_2),
       .op_in      (op_in_0_2),
       .pivot_in   (pivot_in_0_2),
       .start_out  (start_out_0_2),
       .swap_out   (swap_out_0_2),
       .data_out   (data_out_0_2),
       .op_out     (op_out_0_2),
       .pivot_out  (pivot_out_0_2),
       .r          (r_0_2)
     );

  // row 0, col 3

     reg start_in_0_3;
     wire start_out_0_3;

     reg swap_in_0_3;
     wire swap_out_0_3;

     reg [1:0] op_in_0_3;
     wire [1:0] op_out_0_3;

     wire r_0_3;

     wire data_in_0_3;
     wire data_out_0_3;

     reg pivot_in_0_3;
     wire pivot_out_0_3;

     assign data_in_0_3 = data_in[DAT_W-4];

     always @(posedge clk) begin
        op_in_0_3 <= op_out_0_2;
        pivot_in_0_3 <= pivot_out_0_2;
        start_in_0_3 <= start_out_0_2;
        swap_in_0_3 <= swap_out_0_2;
     end
  
     processor_AB AB_0_3 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_3),
       .start_in   (start_in_0_3),
       .swap_in    (swap_in_0_3),
       .op_in      (op_in_0_3),
       .pivot_in   (pivot_in_0_3),
       .start_out  (start_out_0_3),
       .swap_out   (swap_out_0_3),
       .data_out   (data_out_0_3),
       .op_out     (op_out_0_3),
       .pivot_out  (pivot_out_0_3),
       .r          (r_0_3)
     );

  // row 0, col 4

     reg start_in_0_4;
     wire start_out_0_4;

     reg swap_in_0_4;
     wire swap_out_0_4;

     reg [1:0] op_in_0_4;
     wire [1:0] op_out_0_4;

     wire r_0_4;

     wire data_in_0_4;
     wire data_out_0_4;

     reg pivot_in_0_4;
     wire pivot_out_0_4;

     assign data_in_0_4 = data_in[DAT_W-5];

     always @(posedge clk) begin
        op_in_0_4 <= op_out_0_3;
        pivot_in_0_4 <= pivot_out_0_3;
        start_in_0_4 <= start_out_0_3;
        swap_in_0_4 <= swap_out_0_3;
     end
  
     processor_AB AB_0_4 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_4),
       .start_in   (start_in_0_4),
       .swap_in    (swap_in_0_4),
       .op_in      (op_in_0_4),
       .pivot_in   (pivot_in_0_4),
       .start_out  (start_out_0_4),
       .swap_out   (swap_out_0_4),
       .data_out   (data_out_0_4),
       .op_out     (op_out_0_4),
       .pivot_out  (pivot_out_0_4),
       .r          (r_0_4)
     );

  // row 0, col 5

     reg start_in_0_5;
     wire start_out_0_5;

     reg swap_in_0_5;
     wire swap_out_0_5;

     reg [1:0] op_in_0_5;
     wire [1:0] op_out_0_5;

     wire r_0_5;

     wire data_in_0_5;
     wire data_out_0_5;

     reg pivot_in_0_5;
     wire pivot_out_0_5;

     assign data_in_0_5 = data_in[DAT_W-6];

     always @(posedge clk) begin
        op_in_0_5 <= op_out_0_4;
        pivot_in_0_5 <= pivot_out_0_4;
        start_in_0_5 <= start_out_0_4;
        swap_in_0_5 <= swap_out_0_4;
     end
  
     processor_AB AB_0_5 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_5),
       .start_in   (start_in_0_5),
       .swap_in    (swap_in_0_5),
       .op_in      (op_in_0_5),
       .pivot_in   (pivot_in_0_5),
       .start_out  (start_out_0_5),
       .swap_out   (swap_out_0_5),
       .data_out   (data_out_0_5),
       .op_out     (op_out_0_5),
       .pivot_out  (pivot_out_0_5),
       .r          (r_0_5)
     );

  // row 0, col 6

     reg start_in_0_6;
     wire start_out_0_6;

     reg swap_in_0_6;
     wire swap_out_0_6;

     reg [1:0] op_in_0_6;
     wire [1:0] op_out_0_6;

     wire r_0_6;

     wire data_in_0_6;
     wire data_out_0_6;

     reg pivot_in_0_6;
     wire pivot_out_0_6;

     assign data_in_0_6 = data_in[DAT_W-7];

     always @(posedge clk) begin
        op_in_0_6 <= op_out_0_5;
        pivot_in_0_6 <= pivot_out_0_5;
        start_in_0_6 <= start_out_0_5;
        swap_in_0_6 <= swap_out_0_5;
     end
  
     processor_AB AB_0_6 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_6),
       .start_in   (start_in_0_6),
       .swap_in    (swap_in_0_6),
       .op_in      (op_in_0_6),
       .pivot_in   (pivot_in_0_6),
       .start_out  (start_out_0_6),
       .swap_out   (swap_out_0_6),
       .data_out   (data_out_0_6),
       .op_out     (op_out_0_6),
       .pivot_out  (pivot_out_0_6),
       .r          (r_0_6)
     );

  // row 0, col 7

     reg start_in_0_7;
     wire start_out_0_7;

     reg swap_in_0_7;
     wire swap_out_0_7;

     reg [1:0] op_in_0_7;
     wire [1:0] op_out_0_7;

     wire r_0_7;

     wire data_in_0_7;
     wire data_out_0_7;

     reg pivot_in_0_7;
     wire pivot_out_0_7;

     assign data_in_0_7 = data_in[DAT_W-8];

     always @(posedge clk) begin
        op_in_0_7 <= op_out_0_6;
        pivot_in_0_7 <= pivot_out_0_6;
        start_in_0_7 <= start_out_0_6;
        swap_in_0_7 <= swap_out_0_6;
     end
  
     processor_AB AB_0_7 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_7),
       .start_in   (start_in_0_7),
       .swap_in    (swap_in_0_7),
       .op_in      (op_in_0_7),
       .pivot_in   (pivot_in_0_7),
       .start_out  (start_out_0_7),
       .swap_out   (swap_out_0_7),
       .data_out   (data_out_0_7),
       .op_out     (op_out_0_7),
       .pivot_out  (pivot_out_0_7),
       .r          (r_0_7)
     );

  // row 0, col 8

     reg start_in_0_8;
     wire start_out_0_8;

     reg swap_in_0_8;
     wire swap_out_0_8;

     reg [1:0] op_in_0_8;
     wire [1:0] op_out_0_8;

     wire r_0_8;

     wire data_in_0_8;
     wire data_out_0_8;

     reg pivot_in_0_8;
     wire pivot_out_0_8;

     assign data_in_0_8 = data_in[DAT_W-9];

     always @(posedge clk) begin
        op_in_0_8 <= op_out_0_7;
        pivot_in_0_8 <= pivot_out_0_7;
        start_in_0_8 <= start_out_0_7;
        swap_in_0_8 <= swap_out_0_7;
     end
  
     processor_AB AB_0_8 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_8),
       .start_in   (start_in_0_8),
       .swap_in    (swap_in_0_8),
       .op_in      (op_in_0_8),
       .pivot_in   (pivot_in_0_8),
       .start_out  (start_out_0_8),
       .swap_out   (swap_out_0_8),
       .data_out   (data_out_0_8),
       .op_out     (op_out_0_8),
       .pivot_out  (pivot_out_0_8),
       .r          (r_0_8)
     );

  // row 0, col 9

     reg start_in_0_9;
     wire start_out_0_9;

     reg swap_in_0_9;
     wire swap_out_0_9;

     reg [1:0] op_in_0_9;
     wire [1:0] op_out_0_9;

     wire r_0_9;

     wire data_in_0_9;
     wire data_out_0_9;

     reg pivot_in_0_9;
     wire pivot_out_0_9;

     assign data_in_0_9 = data_in[DAT_W-10];

     always @(posedge clk) begin
        op_in_0_9 <= op_out_0_8;
        pivot_in_0_9 <= pivot_out_0_8;
        start_in_0_9 <= start_out_0_8;
        swap_in_0_9 <= swap_out_0_8;
     end
  
     processor_AB AB_0_9 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_9),
       .start_in   (start_in_0_9),
       .swap_in    (swap_in_0_9),
       .op_in      (op_in_0_9),
       .pivot_in   (pivot_in_0_9),
       .start_out  (start_out_0_9),
       .swap_out   (swap_out_0_9),
       .data_out   (data_out_0_9),
       .op_out     (op_out_0_9),
       .pivot_out  (pivot_out_0_9),
       .r          (r_0_9)
     );

  // row 0, col 10

     reg start_in_0_10;
     wire start_out_0_10;

     reg swap_in_0_10;
     wire swap_out_0_10;

     reg [1:0] op_in_0_10;
     wire [1:0] op_out_0_10;

     wire r_0_10;

     wire data_in_0_10;
     wire data_out_0_10;

     reg pivot_in_0_10;
     wire pivot_out_0_10;

     assign data_in_0_10 = data_in[DAT_W-11];

     always @(posedge clk) begin
        op_in_0_10 <= op_out_0_9;
        pivot_in_0_10 <= pivot_out_0_9;
        start_in_0_10 <= start_out_0_9;
        swap_in_0_10 <= swap_out_0_9;
     end
  
     processor_AB AB_0_10 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_10),
       .start_in   (start_in_0_10),
       .swap_in    (swap_in_0_10),
       .op_in      (op_in_0_10),
       .pivot_in   (pivot_in_0_10),
       .start_out  (start_out_0_10),
       .swap_out   (swap_out_0_10),
       .data_out   (data_out_0_10),
       .op_out     (op_out_0_10),
       .pivot_out  (pivot_out_0_10),
       .r          (r_0_10)
     );

  // row 0, col 11

     reg start_in_0_11;
     wire start_out_0_11;

     reg swap_in_0_11;
     wire swap_out_0_11;

     reg [1:0] op_in_0_11;
     wire [1:0] op_out_0_11;

     wire r_0_11;

     wire data_in_0_11;
     wire data_out_0_11;

     reg pivot_in_0_11;
     wire pivot_out_0_11;

     assign data_in_0_11 = data_in[DAT_W-12];

     always @(posedge clk) begin
        op_in_0_11 <= op_out_0_10;
        pivot_in_0_11 <= pivot_out_0_10;
        start_in_0_11 <= start_out_0_10;
        swap_in_0_11 <= swap_out_0_10;
     end
  
     processor_AB AB_0_11 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_11),
       .start_in   (start_in_0_11),
       .swap_in    (swap_in_0_11),
       .op_in      (op_in_0_11),
       .pivot_in   (pivot_in_0_11),
       .start_out  (start_out_0_11),
       .swap_out   (swap_out_0_11),
       .data_out   (data_out_0_11),
       .op_out     (op_out_0_11),
       .pivot_out  (pivot_out_0_11),
       .r          (r_0_11)
     );

  // row 0, col 12

     reg start_in_0_12;
     wire start_out_0_12;

     reg swap_in_0_12;
     wire swap_out_0_12;

     reg [1:0] op_in_0_12;
     wire [1:0] op_out_0_12;

     wire r_0_12;

     wire data_in_0_12;
     wire data_out_0_12;

     reg pivot_in_0_12;
     wire pivot_out_0_12;

     assign data_in_0_12 = data_in[DAT_W-13];

     always @(posedge clk) begin
        op_in_0_12 <= op_out_0_11;
        pivot_in_0_12 <= pivot_out_0_11;
        start_in_0_12 <= start_out_0_11;
        swap_in_0_12 <= swap_out_0_11;
     end
  
     processor_AB AB_0_12 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_12),
       .start_in   (start_in_0_12),
       .swap_in    (swap_in_0_12),
       .op_in      (op_in_0_12),
       .pivot_in   (pivot_in_0_12),
       .start_out  (start_out_0_12),
       .swap_out   (swap_out_0_12),
       .data_out   (data_out_0_12),
       .op_out     (op_out_0_12),
       .pivot_out  (pivot_out_0_12),
       .r          (r_0_12)
     );

  // row 0, col 13

     reg start_in_0_13;
     wire start_out_0_13;

     reg swap_in_0_13;
     wire swap_out_0_13;

     reg [1:0] op_in_0_13;
     wire [1:0] op_out_0_13;

     wire r_0_13;

     wire data_in_0_13;
     wire data_out_0_13;

     reg pivot_in_0_13;
     wire pivot_out_0_13;

     assign data_in_0_13 = data_in[DAT_W-14];

     always @(posedge clk) begin
        op_in_0_13 <= op_out_0_12;
        pivot_in_0_13 <= pivot_out_0_12;
        start_in_0_13 <= start_out_0_12;
        swap_in_0_13 <= swap_out_0_12;
     end
  
     processor_AB AB_0_13 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_13),
       .start_in   (start_in_0_13),
       .swap_in    (swap_in_0_13),
       .op_in      (op_in_0_13),
       .pivot_in   (pivot_in_0_13),
       .start_out  (start_out_0_13),
       .swap_out   (swap_out_0_13),
       .data_out   (data_out_0_13),
       .op_out     (op_out_0_13),
       .pivot_out  (pivot_out_0_13),
       .r          (r_0_13)
     );

  // row 0, col 14

     reg start_in_0_14;
     wire start_out_0_14;

     reg swap_in_0_14;
     wire swap_out_0_14;

     reg [1:0] op_in_0_14;
     wire [1:0] op_out_0_14;

     wire r_0_14;

     wire data_in_0_14;
     wire data_out_0_14;

     reg pivot_in_0_14;
     wire pivot_out_0_14;

     assign data_in_0_14 = data_in[DAT_W-15];

     always @(posedge clk) begin
        op_in_0_14 <= op_out_0_13;
        pivot_in_0_14 <= pivot_out_0_13;
        start_in_0_14 <= start_out_0_13;
        swap_in_0_14 <= swap_out_0_13;
     end
  
     processor_AB AB_0_14 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_14),
       .start_in   (start_in_0_14),
       .swap_in    (swap_in_0_14),
       .op_in      (op_in_0_14),
       .pivot_in   (pivot_in_0_14),
       .start_out  (start_out_0_14),
       .swap_out   (swap_out_0_14),
       .data_out   (data_out_0_14),
       .op_out     (op_out_0_14),
       .pivot_out  (pivot_out_0_14),
       .r          (r_0_14)
     );

  // row 0, col 15

     reg start_in_0_15;
     wire start_out_0_15;

     reg swap_in_0_15;
     wire swap_out_0_15;

     reg [1:0] op_in_0_15;
     wire [1:0] op_out_0_15;

     wire r_0_15;

     wire data_in_0_15;
     wire data_out_0_15;

     reg pivot_in_0_15;
     wire pivot_out_0_15;

     assign data_in_0_15 = data_in[DAT_W-16];

     always @(posedge clk) begin
        op_in_0_15 <= op_out_0_14;
        pivot_in_0_15 <= pivot_out_0_14;
        start_in_0_15 <= start_out_0_14;
        swap_in_0_15 <= swap_out_0_14;
     end
  
     processor_AB AB_0_15 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_15),
       .start_in   (start_in_0_15),
       .swap_in    (swap_in_0_15),
       .op_in      (op_in_0_15),
       .pivot_in   (pivot_in_0_15),
       .start_out  (start_out_0_15),
       .swap_out   (swap_out_0_15),
       .data_out   (data_out_0_15),
       .op_out     (op_out_0_15),
       .pivot_out  (pivot_out_0_15),
       .r          (r_0_15)
     );

  // row 0, col 16

     reg start_in_0_16;
     wire start_out_0_16;

     reg swap_in_0_16;
     wire swap_out_0_16;

     reg [1:0] op_in_0_16;
     wire [1:0] op_out_0_16;

     wire r_0_16;

     wire data_in_0_16;
     wire data_out_0_16;

     reg pivot_in_0_16;
     wire pivot_out_0_16;

     assign data_in_0_16 = data_in[DAT_W-17];

     always @(posedge clk) begin
        op_in_0_16 <= op_out_0_15;
        pivot_in_0_16 <= pivot_out_0_15;
        start_in_0_16 <= start_out_0_15;
        swap_in_0_16 <= swap_out_0_15;
     end
  
     processor_AB AB_0_16 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_16),
       .start_in   (start_in_0_16),
       .swap_in    (swap_in_0_16),
       .op_in      (op_in_0_16),
       .pivot_in   (pivot_in_0_16),
       .start_out  (start_out_0_16),
       .swap_out   (swap_out_0_16),
       .data_out   (data_out_0_16),
       .op_out     (op_out_0_16),
       .pivot_out  (pivot_out_0_16),
       .r          (r_0_16)
     );

  // row 0, col 17

     reg start_in_0_17;
     wire start_out_0_17;

     reg swap_in_0_17;
     wire swap_out_0_17;

     reg [1:0] op_in_0_17;
     wire [1:0] op_out_0_17;

     wire r_0_17;

     wire data_in_0_17;
     wire data_out_0_17;

     reg pivot_in_0_17;
     wire pivot_out_0_17;

     assign data_in_0_17 = data_in[DAT_W-18];

     always @(posedge clk) begin
        op_in_0_17 <= op_out_0_16;
        pivot_in_0_17 <= pivot_out_0_16;
        start_in_0_17 <= start_out_0_16;
        swap_in_0_17 <= swap_out_0_16;
     end
  
     processor_AB AB_0_17 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_17),
       .start_in   (start_in_0_17),
       .swap_in    (swap_in_0_17),
       .op_in      (op_in_0_17),
       .pivot_in   (pivot_in_0_17),
       .start_out  (start_out_0_17),
       .swap_out   (swap_out_0_17),
       .data_out   (data_out_0_17),
       .op_out     (op_out_0_17),
       .pivot_out  (pivot_out_0_17),
       .r          (r_0_17)
     );

  // row 0, col 18

     reg start_in_0_18;
     wire start_out_0_18;

     reg swap_in_0_18;
     wire swap_out_0_18;

     reg [1:0] op_in_0_18;
     wire [1:0] op_out_0_18;

     wire r_0_18;

     wire data_in_0_18;
     wire data_out_0_18;

     reg pivot_in_0_18;
     wire pivot_out_0_18;

     assign data_in_0_18 = data_in[DAT_W-19];

     always @(posedge clk) begin
        op_in_0_18 <= op_out_0_17;
        pivot_in_0_18 <= pivot_out_0_17;
        start_in_0_18 <= start_out_0_17;
        swap_in_0_18 <= swap_out_0_17;
     end
  
     processor_AB AB_0_18 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_18),
       .start_in   (start_in_0_18),
       .swap_in    (swap_in_0_18),
       .op_in      (op_in_0_18),
       .pivot_in   (pivot_in_0_18),
       .start_out  (start_out_0_18),
       .swap_out   (swap_out_0_18),
       .data_out   (data_out_0_18),
       .op_out     (op_out_0_18),
       .pivot_out  (pivot_out_0_18),
       .r          (r_0_18)
     );

  // row 0, col 19

     reg start_in_0_19;
     wire start_out_0_19;

     reg swap_in_0_19;
     wire swap_out_0_19;

     reg [1:0] op_in_0_19;
     wire [1:0] op_out_0_19;

     wire r_0_19;

     wire data_in_0_19;
     wire data_out_0_19;

     reg pivot_in_0_19;
     wire pivot_out_0_19;

     assign data_in_0_19 = data_in[DAT_W-20];

     always @(posedge clk) begin
        op_in_0_19 <= op_out_0_18;
        pivot_in_0_19 <= pivot_out_0_18;
        start_in_0_19 <= start_out_0_18;
        swap_in_0_19 <= swap_out_0_18;
     end
  
     processor_AB AB_0_19 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_19),
       .start_in   (start_in_0_19),
       .swap_in    (swap_in_0_19),
       .op_in      (op_in_0_19),
       .pivot_in   (pivot_in_0_19),
       .start_out  (start_out_0_19),
       .swap_out   (swap_out_0_19),
       .data_out   (data_out_0_19),
       .op_out     (op_out_0_19),
       .pivot_out  (pivot_out_0_19),
       .r          (r_0_19)
     );

  // row 0, col 20

     reg start_in_0_20;
     wire start_out_0_20;

     reg swap_in_0_20;
     wire swap_out_0_20;

     reg [1:0] op_in_0_20;
     wire [1:0] op_out_0_20;

     wire r_0_20;

     wire data_in_0_20;
     wire data_out_0_20;

     reg pivot_in_0_20;
     wire pivot_out_0_20;

     assign data_in_0_20 = data_in[DAT_W-21];

     always @(posedge clk) begin
        op_in_0_20 <= op_out_0_19;
        pivot_in_0_20 <= pivot_out_0_19;
        start_in_0_20 <= start_out_0_19;
        swap_in_0_20 <= swap_out_0_19;
     end
  
     processor_AB AB_0_20 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_20),
       .start_in   (start_in_0_20),
       .swap_in    (swap_in_0_20),
       .op_in      (op_in_0_20),
       .pivot_in   (pivot_in_0_20),
       .start_out  (start_out_0_20),
       .swap_out   (swap_out_0_20),
       .data_out   (data_out_0_20),
       .op_out     (op_out_0_20),
       .pivot_out  (pivot_out_0_20),
       .r          (r_0_20)
     );

  // row 0, col 21

     reg start_in_0_21;
     wire start_out_0_21;

     reg swap_in_0_21;
     wire swap_out_0_21;

     reg [1:0] op_in_0_21;
     wire [1:0] op_out_0_21;

     wire r_0_21;

     wire data_in_0_21;
     wire data_out_0_21;

     reg pivot_in_0_21;
     wire pivot_out_0_21;

     assign data_in_0_21 = data_in[DAT_W-22];

     always @(posedge clk) begin
        op_in_0_21 <= op_out_0_20;
        pivot_in_0_21 <= pivot_out_0_20;
        start_in_0_21 <= start_out_0_20;
        swap_in_0_21 <= swap_out_0_20;
     end
  
     processor_AB AB_0_21 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_21),
       .start_in   (start_in_0_21),
       .swap_in    (swap_in_0_21),
       .op_in      (op_in_0_21),
       .pivot_in   (pivot_in_0_21),
       .start_out  (start_out_0_21),
       .swap_out   (swap_out_0_21),
       .data_out   (data_out_0_21),
       .op_out     (op_out_0_21),
       .pivot_out  (pivot_out_0_21),
       .r          (r_0_21)
     );

  // row 0, col 22

     reg start_in_0_22;
     wire start_out_0_22;

     reg swap_in_0_22;
     wire swap_out_0_22;

     reg [1:0] op_in_0_22;
     wire [1:0] op_out_0_22;

     wire r_0_22;

     wire data_in_0_22;
     wire data_out_0_22;

     reg pivot_in_0_22;
     wire pivot_out_0_22;

     assign data_in_0_22 = data_in[DAT_W-23];

     always @(posedge clk) begin
        op_in_0_22 <= op_out_0_21;
        pivot_in_0_22 <= pivot_out_0_21;
        start_in_0_22 <= start_out_0_21;
        swap_in_0_22 <= swap_out_0_21;
     end
  
     processor_AB AB_0_22 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_22),
       .start_in   (start_in_0_22),
       .swap_in    (swap_in_0_22),
       .op_in      (op_in_0_22),
       .pivot_in   (pivot_in_0_22),
       .start_out  (start_out_0_22),
       .swap_out   (swap_out_0_22),
       .data_out   (data_out_0_22),
       .op_out     (op_out_0_22),
       .pivot_out  (pivot_out_0_22),
       .r          (r_0_22)
     );

  // row 0, col 23

     reg start_in_0_23;
     wire start_out_0_23;

     reg swap_in_0_23;
     wire swap_out_0_23;

     reg [1:0] op_in_0_23;
     wire [1:0] op_out_0_23;

     wire r_0_23;

     wire data_in_0_23;
     wire data_out_0_23;

     reg pivot_in_0_23;
     wire pivot_out_0_23;

     assign data_in_0_23 = data_in[DAT_W-24];

     always @(posedge clk) begin
        op_in_0_23 <= op_out_0_22;
        pivot_in_0_23 <= pivot_out_0_22;
        start_in_0_23 <= start_out_0_22;
        swap_in_0_23 <= swap_out_0_22;
     end
  
     processor_AB AB_0_23 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_23),
       .start_in   (start_in_0_23),
       .swap_in    (swap_in_0_23),
       .op_in      (op_in_0_23),
       .pivot_in   (pivot_in_0_23),
       .start_out  (start_out_0_23),
       .swap_out   (swap_out_0_23),
       .data_out   (data_out_0_23),
       .op_out     (op_out_0_23),
       .pivot_out  (pivot_out_0_23),
       .r          (r_0_23)
     );

  // row 0, col 24

     reg start_in_0_24;
     wire start_out_0_24;

     reg swap_in_0_24;
     wire swap_out_0_24;

     reg [1:0] op_in_0_24;
     wire [1:0] op_out_0_24;

     wire r_0_24;

     wire data_in_0_24;
     wire data_out_0_24;

     reg pivot_in_0_24;
     wire pivot_out_0_24;

     assign data_in_0_24 = data_in[DAT_W-25];

     always @(posedge clk) begin
        op_in_0_24 <= op_out_0_23;
        pivot_in_0_24 <= pivot_out_0_23;
        start_in_0_24 <= start_out_0_23;
        swap_in_0_24 <= swap_out_0_23;
     end
  
     processor_AB AB_0_24 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_24),
       .start_in   (start_in_0_24),
       .swap_in    (swap_in_0_24),
       .op_in      (op_in_0_24),
       .pivot_in   (pivot_in_0_24),
       .start_out  (start_out_0_24),
       .swap_out   (swap_out_0_24),
       .data_out   (data_out_0_24),
       .op_out     (op_out_0_24),
       .pivot_out  (pivot_out_0_24),
       .r          (r_0_24)
     );

  // row 0, col 25

     reg start_in_0_25;
     wire start_out_0_25;

     reg swap_in_0_25;
     wire swap_out_0_25;

     reg [1:0] op_in_0_25;
     wire [1:0] op_out_0_25;

     wire r_0_25;

     wire data_in_0_25;
     wire data_out_0_25;

     reg pivot_in_0_25;
     wire pivot_out_0_25;

     assign data_in_0_25 = data_in[DAT_W-26];

     always @(posedge clk) begin
        op_in_0_25 <= op_out_0_24;
        pivot_in_0_25 <= pivot_out_0_24;
        start_in_0_25 <= start_out_0_24;
        swap_in_0_25 <= swap_out_0_24;
     end
  
     processor_AB AB_0_25 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_25),
       .start_in   (start_in_0_25),
       .swap_in    (swap_in_0_25),
       .op_in      (op_in_0_25),
       .pivot_in   (pivot_in_0_25),
       .start_out  (start_out_0_25),
       .swap_out   (swap_out_0_25),
       .data_out   (data_out_0_25),
       .op_out     (op_out_0_25),
       .pivot_out  (pivot_out_0_25),
       .r          (r_0_25)
     );

  // row 0, col 26

     reg start_in_0_26;
     wire start_out_0_26;

     reg swap_in_0_26;
     wire swap_out_0_26;

     reg [1:0] op_in_0_26;
     wire [1:0] op_out_0_26;

     wire r_0_26;

     wire data_in_0_26;
     wire data_out_0_26;

     reg pivot_in_0_26;
     wire pivot_out_0_26;

     assign data_in_0_26 = data_in[DAT_W-27];

     always @(posedge clk) begin
        op_in_0_26 <= op_out_0_25;
        pivot_in_0_26 <= pivot_out_0_25;
        start_in_0_26 <= start_out_0_25;
        swap_in_0_26 <= swap_out_0_25;
     end
  
     processor_AB AB_0_26 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_26),
       .start_in   (start_in_0_26),
       .swap_in    (swap_in_0_26),
       .op_in      (op_in_0_26),
       .pivot_in   (pivot_in_0_26),
       .start_out  (start_out_0_26),
       .swap_out   (swap_out_0_26),
       .data_out   (data_out_0_26),
       .op_out     (op_out_0_26),
       .pivot_out  (pivot_out_0_26),
       .r          (r_0_26)
     );

  // row 0, col 27

     reg start_in_0_27;
     wire start_out_0_27;

     reg swap_in_0_27;
     wire swap_out_0_27;

     reg [1:0] op_in_0_27;
     wire [1:0] op_out_0_27;

     wire r_0_27;

     wire data_in_0_27;
     wire data_out_0_27;

     reg pivot_in_0_27;
     wire pivot_out_0_27;

     assign data_in_0_27 = data_in[DAT_W-28];

     always @(posedge clk) begin
        op_in_0_27 <= op_out_0_26;
        pivot_in_0_27 <= pivot_out_0_26;
        start_in_0_27 <= start_out_0_26;
        swap_in_0_27 <= swap_out_0_26;
     end
  
     processor_AB AB_0_27 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_27),
       .start_in   (start_in_0_27),
       .swap_in    (swap_in_0_27),
       .op_in      (op_in_0_27),
       .pivot_in   (pivot_in_0_27),
       .start_out  (start_out_0_27),
       .swap_out   (swap_out_0_27),
       .data_out   (data_out_0_27),
       .op_out     (op_out_0_27),
       .pivot_out  (pivot_out_0_27),
       .r          (r_0_27)
     );

  // row 0, col 28

     reg start_in_0_28;
     wire start_out_0_28;

     reg swap_in_0_28;
     wire swap_out_0_28;

     reg [1:0] op_in_0_28;
     wire [1:0] op_out_0_28;

     wire r_0_28;

     wire data_in_0_28;
     wire data_out_0_28;

     reg pivot_in_0_28;
     wire pivot_out_0_28;

     assign data_in_0_28 = data_in[DAT_W-29];

     always @(posedge clk) begin
        op_in_0_28 <= op_out_0_27;
        pivot_in_0_28 <= pivot_out_0_27;
        start_in_0_28 <= start_out_0_27;
        swap_in_0_28 <= swap_out_0_27;
     end
  
     processor_AB AB_0_28 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_28),
       .start_in   (start_in_0_28),
       .swap_in    (swap_in_0_28),
       .op_in      (op_in_0_28),
       .pivot_in   (pivot_in_0_28),
       .start_out  (start_out_0_28),
       .swap_out   (swap_out_0_28),
       .data_out   (data_out_0_28),
       .op_out     (op_out_0_28),
       .pivot_out  (pivot_out_0_28),
       .r          (r_0_28)
     );

  // row 0, col 29

     reg start_in_0_29;
     wire start_out_0_29;

     reg swap_in_0_29;
     wire swap_out_0_29;

     reg [1:0] op_in_0_29;
     wire [1:0] op_out_0_29;

     wire r_0_29;

     wire data_in_0_29;
     wire data_out_0_29;

     reg pivot_in_0_29;
     wire pivot_out_0_29;

     assign data_in_0_29 = data_in[DAT_W-30];

     always @(posedge clk) begin
        op_in_0_29 <= op_out_0_28;
        pivot_in_0_29 <= pivot_out_0_28;
        start_in_0_29 <= start_out_0_28;
        swap_in_0_29 <= swap_out_0_28;
     end
  
     processor_AB AB_0_29 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_29),
       .start_in   (start_in_0_29),
       .swap_in    (swap_in_0_29),
       .op_in      (op_in_0_29),
       .pivot_in   (pivot_in_0_29),
       .start_out  (start_out_0_29),
       .swap_out   (swap_out_0_29),
       .data_out   (data_out_0_29),
       .op_out     (op_out_0_29),
       .pivot_out  (pivot_out_0_29),
       .r          (r_0_29)
     );

  // row 0, col 30

     reg start_in_0_30;
     wire start_out_0_30;

     reg swap_in_0_30;
     wire swap_out_0_30;

     reg [1:0] op_in_0_30;
     wire [1:0] op_out_0_30;

     wire r_0_30;

     wire data_in_0_30;
     wire data_out_0_30;

     reg pivot_in_0_30;
     wire pivot_out_0_30;

     assign data_in_0_30 = data_in[DAT_W-31];

     always @(posedge clk) begin
        op_in_0_30 <= op_out_0_29;
        pivot_in_0_30 <= pivot_out_0_29;
        start_in_0_30 <= start_out_0_29;
        swap_in_0_30 <= swap_out_0_29;
     end
  
     processor_AB AB_0_30 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_30),
       .start_in   (start_in_0_30),
       .swap_in    (swap_in_0_30),
       .op_in      (op_in_0_30),
       .pivot_in   (pivot_in_0_30),
       .start_out  (start_out_0_30),
       .swap_out   (swap_out_0_30),
       .data_out   (data_out_0_30),
       .op_out     (op_out_0_30),
       .pivot_out  (pivot_out_0_30),
       .r          (r_0_30)
     );

  // row 0, col 31

     reg start_in_0_31;
     wire start_out_0_31;

     reg swap_in_0_31;
     wire swap_out_0_31;

     reg [1:0] op_in_0_31;
     wire [1:0] op_out_0_31;

     wire r_0_31;

     wire data_in_0_31;
     wire data_out_0_31;

     reg pivot_in_0_31;
     wire pivot_out_0_31;

     assign data_in_0_31 = data_in[DAT_W-32];

     always @(posedge clk) begin
        op_in_0_31 <= op_out_0_30;
        pivot_in_0_31 <= pivot_out_0_30;
        start_in_0_31 <= start_out_0_30;
        swap_in_0_31 <= swap_out_0_30;
     end
  
     processor_AB AB_0_31 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_31),
       .start_in   (start_in_0_31),
       .swap_in    (swap_in_0_31),
       .op_in      (op_in_0_31),
       .pivot_in   (pivot_in_0_31),
       .start_out  (start_out_0_31),
       .swap_out   (swap_out_0_31),
       .data_out   (data_out_0_31),
       .op_out     (op_out_0_31),
       .pivot_out  (pivot_out_0_31),
       .r          (r_0_31)
     );

  // row 0, col 32

     reg start_in_0_32;
     wire start_out_0_32;

     reg swap_in_0_32;
     wire swap_out_0_32;

     reg [1:0] op_in_0_32;
     wire [1:0] op_out_0_32;

     wire r_0_32;

     wire data_in_0_32;
     wire data_out_0_32;

     reg pivot_in_0_32;
     wire pivot_out_0_32;

     assign data_in_0_32 = data_in[DAT_W-33];

     always @(posedge clk) begin
        op_in_0_32 <= op_out_0_31;
        pivot_in_0_32 <= pivot_out_0_31;
        start_in_0_32 <= start_out_0_31;
        swap_in_0_32 <= swap_out_0_31;
     end
  
     processor_AB AB_0_32 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_32),
       .start_in   (start_in_0_32),
       .swap_in    (swap_in_0_32),
       .op_in      (op_in_0_32),
       .pivot_in   (pivot_in_0_32),
       .start_out  (start_out_0_32),
       .swap_out   (swap_out_0_32),
       .data_out   (data_out_0_32),
       .op_out     (op_out_0_32),
       .pivot_out  (pivot_out_0_32),
       .r          (r_0_32)
     );

  // row 0, col 33

     reg start_in_0_33;
     wire start_out_0_33;

     reg swap_in_0_33;
     wire swap_out_0_33;

     reg [1:0] op_in_0_33;
     wire [1:0] op_out_0_33;

     wire r_0_33;

     wire data_in_0_33;
     wire data_out_0_33;

     reg pivot_in_0_33;
     wire pivot_out_0_33;

     assign data_in_0_33 = data_in[DAT_W-34];

     always @(posedge clk) begin
        op_in_0_33 <= op_out_0_32;
        pivot_in_0_33 <= pivot_out_0_32;
        start_in_0_33 <= start_out_0_32;
        swap_in_0_33 <= swap_out_0_32;
     end
  
     processor_AB AB_0_33 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_33),
       .start_in   (start_in_0_33),
       .swap_in    (swap_in_0_33),
       .op_in      (op_in_0_33),
       .pivot_in   (pivot_in_0_33),
       .start_out  (start_out_0_33),
       .swap_out   (swap_out_0_33),
       .data_out   (data_out_0_33),
       .op_out     (op_out_0_33),
       .pivot_out  (pivot_out_0_33),
       .r          (r_0_33)
     );

  // row 0, col 34

     reg start_in_0_34;
     wire start_out_0_34;

     reg swap_in_0_34;
     wire swap_out_0_34;

     reg [1:0] op_in_0_34;
     wire [1:0] op_out_0_34;

     wire r_0_34;

     wire data_in_0_34;
     wire data_out_0_34;

     reg pivot_in_0_34;
     wire pivot_out_0_34;

     assign data_in_0_34 = data_in[DAT_W-35];

     always @(posedge clk) begin
        op_in_0_34 <= op_out_0_33;
        pivot_in_0_34 <= pivot_out_0_33;
        start_in_0_34 <= start_out_0_33;
        swap_in_0_34 <= swap_out_0_33;
     end
  
     processor_AB AB_0_34 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_34),
       .start_in   (start_in_0_34),
       .swap_in    (swap_in_0_34),
       .op_in      (op_in_0_34),
       .pivot_in   (pivot_in_0_34),
       .start_out  (start_out_0_34),
       .swap_out   (swap_out_0_34),
       .data_out   (data_out_0_34),
       .op_out     (op_out_0_34),
       .pivot_out  (pivot_out_0_34),
       .r          (r_0_34)
     );

  // row 0, col 35

     reg start_in_0_35;
     wire start_out_0_35;

     reg swap_in_0_35;
     wire swap_out_0_35;

     reg [1:0] op_in_0_35;
     wire [1:0] op_out_0_35;

     wire r_0_35;

     wire data_in_0_35;
     wire data_out_0_35;

     reg pivot_in_0_35;
     wire pivot_out_0_35;

     assign data_in_0_35 = data_in[DAT_W-36];

     always @(posedge clk) begin
        op_in_0_35 <= op_out_0_34;
        pivot_in_0_35 <= pivot_out_0_34;
        start_in_0_35 <= start_out_0_34;
        swap_in_0_35 <= swap_out_0_34;
     end
  
     processor_AB AB_0_35 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_35),
       .start_in   (start_in_0_35),
       .swap_in    (swap_in_0_35),
       .op_in      (op_in_0_35),
       .pivot_in   (pivot_in_0_35),
       .start_out  (start_out_0_35),
       .swap_out   (swap_out_0_35),
       .data_out   (data_out_0_35),
       .op_out     (op_out_0_35),
       .pivot_out  (pivot_out_0_35),
       .r          (r_0_35)
     );

  // row 0, col 36

     reg start_in_0_36;
     wire start_out_0_36;

     reg swap_in_0_36;
     wire swap_out_0_36;

     reg [1:0] op_in_0_36;
     wire [1:0] op_out_0_36;

     wire r_0_36;

     wire data_in_0_36;
     wire data_out_0_36;

     reg pivot_in_0_36;
     wire pivot_out_0_36;

     assign data_in_0_36 = data_in[DAT_W-37];

     always @(posedge clk) begin
        op_in_0_36 <= op_out_0_35;
        pivot_in_0_36 <= pivot_out_0_35;
        start_in_0_36 <= start_out_0_35;
        swap_in_0_36 <= swap_out_0_35;
     end
  
     processor_AB AB_0_36 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_36),
       .start_in   (start_in_0_36),
       .swap_in    (swap_in_0_36),
       .op_in      (op_in_0_36),
       .pivot_in   (pivot_in_0_36),
       .start_out  (start_out_0_36),
       .swap_out   (swap_out_0_36),
       .data_out   (data_out_0_36),
       .op_out     (op_out_0_36),
       .pivot_out  (pivot_out_0_36),
       .r          (r_0_36)
     );

  // row 0, col 37

     reg start_in_0_37;
     wire start_out_0_37;

     reg swap_in_0_37;
     wire swap_out_0_37;

     reg [1:0] op_in_0_37;
     wire [1:0] op_out_0_37;

     wire r_0_37;

     wire data_in_0_37;
     wire data_out_0_37;

     reg pivot_in_0_37;
     wire pivot_out_0_37;

     assign data_in_0_37 = data_in[DAT_W-38];

     always @(posedge clk) begin
        op_in_0_37 <= op_out_0_36;
        pivot_in_0_37 <= pivot_out_0_36;
        start_in_0_37 <= start_out_0_36;
        swap_in_0_37 <= swap_out_0_36;
     end
  
     processor_AB AB_0_37 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_37),
       .start_in   (start_in_0_37),
       .swap_in    (swap_in_0_37),
       .op_in      (op_in_0_37),
       .pivot_in   (pivot_in_0_37),
       .start_out  (start_out_0_37),
       .swap_out   (swap_out_0_37),
       .data_out   (data_out_0_37),
       .op_out     (op_out_0_37),
       .pivot_out  (pivot_out_0_37),
       .r          (r_0_37)
     );

  // row 0, col 38

     reg start_in_0_38;
     wire start_out_0_38;

     reg swap_in_0_38;
     wire swap_out_0_38;

     reg [1:0] op_in_0_38;
     wire [1:0] op_out_0_38;

     wire r_0_38;

     wire data_in_0_38;
     wire data_out_0_38;

     reg pivot_in_0_38;
     wire pivot_out_0_38;

     assign data_in_0_38 = data_in[DAT_W-39];

     always @(posedge clk) begin
        op_in_0_38 <= op_out_0_37;
        pivot_in_0_38 <= pivot_out_0_37;
        start_in_0_38 <= start_out_0_37;
        swap_in_0_38 <= swap_out_0_37;
     end
  
     processor_AB AB_0_38 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_38),
       .start_in   (start_in_0_38),
       .swap_in    (swap_in_0_38),
       .op_in      (op_in_0_38),
       .pivot_in   (pivot_in_0_38),
       .start_out  (start_out_0_38),
       .swap_out   (swap_out_0_38),
       .data_out   (data_out_0_38),
       .op_out     (op_out_0_38),
       .pivot_out  (pivot_out_0_38),
       .r          (r_0_38)
     );

  // row 0, col 39

     reg start_in_0_39;
     wire start_out_0_39;

     reg swap_in_0_39;
     wire swap_out_0_39;

     reg [1:0] op_in_0_39;
     wire [1:0] op_out_0_39;

     wire r_0_39;

     wire data_in_0_39;
     wire data_out_0_39;

     reg pivot_in_0_39;
     wire pivot_out_0_39;

     assign data_in_0_39 = data_in[DAT_W-40];

     always @(posedge clk) begin
        op_in_0_39 <= op_out_0_38;
        pivot_in_0_39 <= pivot_out_0_38;
        start_in_0_39 <= start_out_0_38;
        swap_in_0_39 <= swap_out_0_38;
     end
  
     processor_AB AB_0_39 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_39),
       .start_in   (start_in_0_39),
       .swap_in    (swap_in_0_39),
       .op_in      (op_in_0_39),
       .pivot_in   (pivot_in_0_39),
       .start_out  (start_out_0_39),
       .swap_out   (swap_out_0_39),
       .data_out   (data_out_0_39),
       .op_out     (op_out_0_39),
       .pivot_out  (pivot_out_0_39),
       .r          (r_0_39)
     );

  // row 0, col 40

     reg start_in_0_40;
     wire start_out_0_40;

     reg swap_in_0_40;
     wire swap_out_0_40;

     reg [1:0] op_in_0_40;
     wire [1:0] op_out_0_40;

     wire r_0_40;

     wire data_in_0_40;
     wire data_out_0_40;

     reg pivot_in_0_40;
     wire pivot_out_0_40;

     assign data_in_0_40 = data_in[DAT_W-41];

     always @(posedge clk) begin
        op_in_0_40 <= op_out_0_39;
        pivot_in_0_40 <= pivot_out_0_39;
        start_in_0_40 <= start_out_0_39;
        swap_in_0_40 <= swap_out_0_39;
     end
  
     processor_AB AB_0_40 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_40),
       .start_in   (start_in_0_40),
       .swap_in    (swap_in_0_40),
       .op_in      (op_in_0_40),
       .pivot_in   (pivot_in_0_40),
       .start_out  (start_out_0_40),
       .swap_out   (swap_out_0_40),
       .data_out   (data_out_0_40),
       .op_out     (op_out_0_40),
       .pivot_out  (pivot_out_0_40),
       .r          (r_0_40)
     );

  // row 0, col 41

     reg start_in_0_41;
     wire start_out_0_41;

     reg swap_in_0_41;
     wire swap_out_0_41;

     reg [1:0] op_in_0_41;
     wire [1:0] op_out_0_41;

     wire r_0_41;

     wire data_in_0_41;
     wire data_out_0_41;

     reg pivot_in_0_41;
     wire pivot_out_0_41;

     assign data_in_0_41 = data_in[DAT_W-42];

     always @(posedge clk) begin
        op_in_0_41 <= op_out_0_40;
        pivot_in_0_41 <= pivot_out_0_40;
        start_in_0_41 <= start_out_0_40;
        swap_in_0_41 <= swap_out_0_40;
     end
  
     processor_AB AB_0_41 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_41),
       .start_in   (start_in_0_41),
       .swap_in    (swap_in_0_41),
       .op_in      (op_in_0_41),
       .pivot_in   (pivot_in_0_41),
       .start_out  (start_out_0_41),
       .swap_out   (swap_out_0_41),
       .data_out   (data_out_0_41),
       .op_out     (op_out_0_41),
       .pivot_out  (pivot_out_0_41),
       .r          (r_0_41)
     );

  // row 0, col 42

     reg start_in_0_42;
     wire start_out_0_42;

     reg swap_in_0_42;
     wire swap_out_0_42;

     reg [1:0] op_in_0_42;
     wire [1:0] op_out_0_42;

     wire r_0_42;

     wire data_in_0_42;
     wire data_out_0_42;

     reg pivot_in_0_42;
     wire pivot_out_0_42;

     assign data_in_0_42 = data_in[DAT_W-43];

     always @(posedge clk) begin
        op_in_0_42 <= op_out_0_41;
        pivot_in_0_42 <= pivot_out_0_41;
        start_in_0_42 <= start_out_0_41;
        swap_in_0_42 <= swap_out_0_41;
     end
  
     processor_AB AB_0_42 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_42),
       .start_in   (start_in_0_42),
       .swap_in    (swap_in_0_42),
       .op_in      (op_in_0_42),
       .pivot_in   (pivot_in_0_42),
       .start_out  (start_out_0_42),
       .swap_out   (swap_out_0_42),
       .data_out   (data_out_0_42),
       .op_out     (op_out_0_42),
       .pivot_out  (pivot_out_0_42),
       .r          (r_0_42)
     );

  // row 0, col 43

     reg start_in_0_43;
     wire start_out_0_43;

     reg swap_in_0_43;
     wire swap_out_0_43;

     reg [1:0] op_in_0_43;
     wire [1:0] op_out_0_43;

     wire r_0_43;

     wire data_in_0_43;
     wire data_out_0_43;

     reg pivot_in_0_43;
     wire pivot_out_0_43;

     assign data_in_0_43 = data_in[DAT_W-44];

     always @(posedge clk) begin
        op_in_0_43 <= op_out_0_42;
        pivot_in_0_43 <= pivot_out_0_42;
        start_in_0_43 <= start_out_0_42;
        swap_in_0_43 <= swap_out_0_42;
     end
  
     processor_AB AB_0_43 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_43),
       .start_in   (start_in_0_43),
       .swap_in    (swap_in_0_43),
       .op_in      (op_in_0_43),
       .pivot_in   (pivot_in_0_43),
       .start_out  (start_out_0_43),
       .swap_out   (swap_out_0_43),
       .data_out   (data_out_0_43),
       .op_out     (op_out_0_43),
       .pivot_out  (pivot_out_0_43),
       .r          (r_0_43)
     );

  // row 0, col 44

     reg start_in_0_44;
     wire start_out_0_44;

     reg swap_in_0_44;
     wire swap_out_0_44;

     reg [1:0] op_in_0_44;
     wire [1:0] op_out_0_44;

     wire r_0_44;

     wire data_in_0_44;
     wire data_out_0_44;

     reg pivot_in_0_44;
     wire pivot_out_0_44;

     assign data_in_0_44 = data_in[DAT_W-45];

     always @(posedge clk) begin
        op_in_0_44 <= op_out_0_43;
        pivot_in_0_44 <= pivot_out_0_43;
        start_in_0_44 <= start_out_0_43;
        swap_in_0_44 <= swap_out_0_43;
     end
  
     processor_AB AB_0_44 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_44),
       .start_in   (start_in_0_44),
       .swap_in    (swap_in_0_44),
       .op_in      (op_in_0_44),
       .pivot_in   (pivot_in_0_44),
       .start_out  (start_out_0_44),
       .swap_out   (swap_out_0_44),
       .data_out   (data_out_0_44),
       .op_out     (op_out_0_44),
       .pivot_out  (pivot_out_0_44),
       .r          (r_0_44)
     );

  // row 0, col 45

     reg start_in_0_45;
     wire start_out_0_45;

     reg swap_in_0_45;
     wire swap_out_0_45;

     reg [1:0] op_in_0_45;
     wire [1:0] op_out_0_45;

     wire r_0_45;

     wire data_in_0_45;
     wire data_out_0_45;

     reg pivot_in_0_45;
     wire pivot_out_0_45;

     assign data_in_0_45 = data_in[DAT_W-46];

     always @(posedge clk) begin
        op_in_0_45 <= op_out_0_44;
        pivot_in_0_45 <= pivot_out_0_44;
        start_in_0_45 <= start_out_0_44;
        swap_in_0_45 <= swap_out_0_44;
     end
  
     processor_AB AB_0_45 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_45),
       .start_in   (start_in_0_45),
       .swap_in    (swap_in_0_45),
       .op_in      (op_in_0_45),
       .pivot_in   (pivot_in_0_45),
       .start_out  (start_out_0_45),
       .swap_out   (swap_out_0_45),
       .data_out   (data_out_0_45),
       .op_out     (op_out_0_45),
       .pivot_out  (pivot_out_0_45),
       .r          (r_0_45)
     );

  // row 0, col 46

     reg start_in_0_46;
     wire start_out_0_46;

     reg swap_in_0_46;
     wire swap_out_0_46;

     reg [1:0] op_in_0_46;
     wire [1:0] op_out_0_46;

     wire r_0_46;

     wire data_in_0_46;
     wire data_out_0_46;

     reg pivot_in_0_46;
     wire pivot_out_0_46;

     assign data_in_0_46 = data_in[DAT_W-47];

     always @(posedge clk) begin
        op_in_0_46 <= op_out_0_45;
        pivot_in_0_46 <= pivot_out_0_45;
        start_in_0_46 <= start_out_0_45;
        swap_in_0_46 <= swap_out_0_45;
     end
  
     processor_AB AB_0_46 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_46),
       .start_in   (start_in_0_46),
       .swap_in    (swap_in_0_46),
       .op_in      (op_in_0_46),
       .pivot_in   (pivot_in_0_46),
       .start_out  (start_out_0_46),
       .swap_out   (swap_out_0_46),
       .data_out   (data_out_0_46),
       .op_out     (op_out_0_46),
       .pivot_out  (pivot_out_0_46),
       .r          (r_0_46)
     );

  // row 0, col 47

     reg start_in_0_47;
     wire start_out_0_47;

     reg swap_in_0_47;
     wire swap_out_0_47;

     reg [1:0] op_in_0_47;
     wire [1:0] op_out_0_47;

     wire r_0_47;

     wire data_in_0_47;
     wire data_out_0_47;

     reg pivot_in_0_47;
     wire pivot_out_0_47;

     assign data_in_0_47 = data_in[DAT_W-48];

     always @(posedge clk) begin
        op_in_0_47 <= op_out_0_46;
        pivot_in_0_47 <= pivot_out_0_46;
        start_in_0_47 <= start_out_0_46;
        swap_in_0_47 <= swap_out_0_46;
     end
  
     processor_AB AB_0_47 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_47),
       .start_in   (start_in_0_47),
       .swap_in    (swap_in_0_47),
       .op_in      (op_in_0_47),
       .pivot_in   (pivot_in_0_47),
       .start_out  (start_out_0_47),
       .swap_out   (swap_out_0_47),
       .data_out   (data_out_0_47),
       .op_out     (op_out_0_47),
       .pivot_out  (pivot_out_0_47),
       .r          (r_0_47)
     );

  // row 0, col 48

     reg start_in_0_48;
     wire start_out_0_48;

     reg swap_in_0_48;
     wire swap_out_0_48;

     reg [1:0] op_in_0_48;
     wire [1:0] op_out_0_48;

     wire r_0_48;

     wire data_in_0_48;
     wire data_out_0_48;

     reg pivot_in_0_48;
     wire pivot_out_0_48;

     assign data_in_0_48 = data_in[DAT_W-49];

     always @(posedge clk) begin
        op_in_0_48 <= op_out_0_47;
        pivot_in_0_48 <= pivot_out_0_47;
        start_in_0_48 <= start_out_0_47;
        swap_in_0_48 <= swap_out_0_47;
     end
  
     processor_AB AB_0_48 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_48),
       .start_in   (start_in_0_48),
       .swap_in    (swap_in_0_48),
       .op_in      (op_in_0_48),
       .pivot_in   (pivot_in_0_48),
       .start_out  (start_out_0_48),
       .swap_out   (swap_out_0_48),
       .data_out   (data_out_0_48),
       .op_out     (op_out_0_48),
       .pivot_out  (pivot_out_0_48),
       .r          (r_0_48)
     );

  // row 0, col 49

     reg start_in_0_49;
     wire start_out_0_49;

     reg swap_in_0_49;
     wire swap_out_0_49;

     reg [1:0] op_in_0_49;
     wire [1:0] op_out_0_49;

     wire r_0_49;

     wire data_in_0_49;
     wire data_out_0_49;

     reg pivot_in_0_49;
     wire pivot_out_0_49;

     assign data_in_0_49 = data_in[DAT_W-50];

     always @(posedge clk) begin
        op_in_0_49 <= op_out_0_48;
        pivot_in_0_49 <= pivot_out_0_48;
        start_in_0_49 <= start_out_0_48;
        swap_in_0_49 <= swap_out_0_48;
     end
  
     processor_AB AB_0_49 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_49),
       .start_in   (start_in_0_49),
       .swap_in    (swap_in_0_49),
       .op_in      (op_in_0_49),
       .pivot_in   (pivot_in_0_49),
       .start_out  (start_out_0_49),
       .swap_out   (swap_out_0_49),
       .data_out   (data_out_0_49),
       .op_out     (op_out_0_49),
       .pivot_out  (pivot_out_0_49),
       .r          (r_0_49)
     );

  // row 0, col 50

     reg start_in_0_50;
     wire start_out_0_50;

     reg swap_in_0_50;
     wire swap_out_0_50;

     reg [1:0] op_in_0_50;
     wire [1:0] op_out_0_50;

     wire r_0_50;

     wire data_in_0_50;
     wire data_out_0_50;

     reg pivot_in_0_50;
     wire pivot_out_0_50;

     assign data_in_0_50 = data_in[DAT_W-51];

     always @(posedge clk) begin
        op_in_0_50 <= op_out_0_49;
        pivot_in_0_50 <= pivot_out_0_49;
        start_in_0_50 <= start_out_0_49;
        swap_in_0_50 <= swap_out_0_49;
     end
  
     processor_AB AB_0_50 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_50),
       .start_in   (start_in_0_50),
       .swap_in    (swap_in_0_50),
       .op_in      (op_in_0_50),
       .pivot_in   (pivot_in_0_50),
       .start_out  (start_out_0_50),
       .swap_out   (swap_out_0_50),
       .data_out   (data_out_0_50),
       .op_out     (op_out_0_50),
       .pivot_out  (pivot_out_0_50),
       .r          (r_0_50)
     );

  // row 0, col 51

     reg start_in_0_51;
     wire start_out_0_51;

     reg swap_in_0_51;
     wire swap_out_0_51;

     reg [1:0] op_in_0_51;
     wire [1:0] op_out_0_51;

     wire r_0_51;

     wire data_in_0_51;
     wire data_out_0_51;

     reg pivot_in_0_51;
     wire pivot_out_0_51;

     assign data_in_0_51 = data_in[DAT_W-52];

     always @(posedge clk) begin
        op_in_0_51 <= op_out_0_50;
        pivot_in_0_51 <= pivot_out_0_50;
        start_in_0_51 <= start_out_0_50;
        swap_in_0_51 <= swap_out_0_50;
     end
  
     processor_AB AB_0_51 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_51),
       .start_in   (start_in_0_51),
       .swap_in    (swap_in_0_51),
       .op_in      (op_in_0_51),
       .pivot_in   (pivot_in_0_51),
       .start_out  (start_out_0_51),
       .swap_out   (swap_out_0_51),
       .data_out   (data_out_0_51),
       .op_out     (op_out_0_51),
       .pivot_out  (pivot_out_0_51),
       .r          (r_0_51)
     );

  // row 0, col 52

     reg start_in_0_52;
     wire start_out_0_52;

     reg swap_in_0_52;
     wire swap_out_0_52;

     reg [1:0] op_in_0_52;
     wire [1:0] op_out_0_52;

     wire r_0_52;

     wire data_in_0_52;
     wire data_out_0_52;

     reg pivot_in_0_52;
     wire pivot_out_0_52;

     assign data_in_0_52 = data_in[DAT_W-53];

     always @(posedge clk) begin
        op_in_0_52 <= op_out_0_51;
        pivot_in_0_52 <= pivot_out_0_51;
        start_in_0_52 <= start_out_0_51;
        swap_in_0_52 <= swap_out_0_51;
     end
  
     processor_AB AB_0_52 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_52),
       .start_in   (start_in_0_52),
       .swap_in    (swap_in_0_52),
       .op_in      (op_in_0_52),
       .pivot_in   (pivot_in_0_52),
       .start_out  (start_out_0_52),
       .swap_out   (swap_out_0_52),
       .data_out   (data_out_0_52),
       .op_out     (op_out_0_52),
       .pivot_out  (pivot_out_0_52),
       .r          (r_0_52)
     );

  // row 0, col 53

     reg start_in_0_53;
     wire start_out_0_53;

     reg swap_in_0_53;
     wire swap_out_0_53;

     reg [1:0] op_in_0_53;
     wire [1:0] op_out_0_53;

     wire r_0_53;

     wire data_in_0_53;
     wire data_out_0_53;

     reg pivot_in_0_53;
     wire pivot_out_0_53;

     assign data_in_0_53 = data_in[DAT_W-54];

     always @(posedge clk) begin
        op_in_0_53 <= op_out_0_52;
        pivot_in_0_53 <= pivot_out_0_52;
        start_in_0_53 <= start_out_0_52;
        swap_in_0_53 <= swap_out_0_52;
     end
  
     processor_AB AB_0_53 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_53),
       .start_in   (start_in_0_53),
       .swap_in    (swap_in_0_53),
       .op_in      (op_in_0_53),
       .pivot_in   (pivot_in_0_53),
       .start_out  (start_out_0_53),
       .swap_out   (swap_out_0_53),
       .data_out   (data_out_0_53),
       .op_out     (op_out_0_53),
       .pivot_out  (pivot_out_0_53),
       .r          (r_0_53)
     );

  // row 0, col 54

     reg start_in_0_54;
     wire start_out_0_54;

     reg swap_in_0_54;
     wire swap_out_0_54;

     reg [1:0] op_in_0_54;
     wire [1:0] op_out_0_54;

     wire r_0_54;

     wire data_in_0_54;
     wire data_out_0_54;

     reg pivot_in_0_54;
     wire pivot_out_0_54;

     assign data_in_0_54 = data_in[DAT_W-55];

     always @(posedge clk) begin
        op_in_0_54 <= op_out_0_53;
        pivot_in_0_54 <= pivot_out_0_53;
        start_in_0_54 <= start_out_0_53;
        swap_in_0_54 <= swap_out_0_53;
     end
  
     processor_AB AB_0_54 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_54),
       .start_in   (start_in_0_54),
       .swap_in    (swap_in_0_54),
       .op_in      (op_in_0_54),
       .pivot_in   (pivot_in_0_54),
       .start_out  (start_out_0_54),
       .swap_out   (swap_out_0_54),
       .data_out   (data_out_0_54),
       .op_out     (op_out_0_54),
       .pivot_out  (pivot_out_0_54),
       .r          (r_0_54)
     );

  // row 0, col 55

     reg start_in_0_55;
     wire start_out_0_55;

     reg swap_in_0_55;
     wire swap_out_0_55;

     reg [1:0] op_in_0_55;
     wire [1:0] op_out_0_55;

     wire r_0_55;

     wire data_in_0_55;
     wire data_out_0_55;

     reg pivot_in_0_55;
     wire pivot_out_0_55;

     assign data_in_0_55 = data_in[DAT_W-56];

     always @(posedge clk) begin
        op_in_0_55 <= op_out_0_54;
        pivot_in_0_55 <= pivot_out_0_54;
        start_in_0_55 <= start_out_0_54;
        swap_in_0_55 <= swap_out_0_54;
     end
  
     processor_AB AB_0_55 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_55),
       .start_in   (start_in_0_55),
       .swap_in    (swap_in_0_55),
       .op_in      (op_in_0_55),
       .pivot_in   (pivot_in_0_55),
       .start_out  (start_out_0_55),
       .swap_out   (swap_out_0_55),
       .data_out   (data_out_0_55),
       .op_out     (op_out_0_55),
       .pivot_out  (pivot_out_0_55),
       .r          (r_0_55)
     );

  // row 0, col 56

     reg start_in_0_56;
     wire start_out_0_56;

     reg swap_in_0_56;
     wire swap_out_0_56;

     reg [1:0] op_in_0_56;
     wire [1:0] op_out_0_56;

     wire r_0_56;

     wire data_in_0_56;
     wire data_out_0_56;

     reg pivot_in_0_56;
     wire pivot_out_0_56;

     assign data_in_0_56 = data_in[DAT_W-57];

     always @(posedge clk) begin
        op_in_0_56 <= op_out_0_55;
        pivot_in_0_56 <= pivot_out_0_55;
        start_in_0_56 <= start_out_0_55;
        swap_in_0_56 <= swap_out_0_55;
     end
  
     processor_AB AB_0_56 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_56),
       .start_in   (start_in_0_56),
       .swap_in    (swap_in_0_56),
       .op_in      (op_in_0_56),
       .pivot_in   (pivot_in_0_56),
       .start_out  (start_out_0_56),
       .swap_out   (swap_out_0_56),
       .data_out   (data_out_0_56),
       .op_out     (op_out_0_56),
       .pivot_out  (pivot_out_0_56),
       .r          (r_0_56)
     );

  // row 0, col 57

     reg start_in_0_57;
     wire start_out_0_57;

     reg swap_in_0_57;
     wire swap_out_0_57;

     reg [1:0] op_in_0_57;
     wire [1:0] op_out_0_57;

     wire r_0_57;

     wire data_in_0_57;
     wire data_out_0_57;

     reg pivot_in_0_57;
     wire pivot_out_0_57;

     assign data_in_0_57 = data_in[DAT_W-58];

     always @(posedge clk) begin
        op_in_0_57 <= op_out_0_56;
        pivot_in_0_57 <= pivot_out_0_56;
        start_in_0_57 <= start_out_0_56;
        swap_in_0_57 <= swap_out_0_56;
     end
  
     processor_AB AB_0_57 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_57),
       .start_in   (start_in_0_57),
       .swap_in    (swap_in_0_57),
       .op_in      (op_in_0_57),
       .pivot_in   (pivot_in_0_57),
       .start_out  (start_out_0_57),
       .swap_out   (swap_out_0_57),
       .data_out   (data_out_0_57),
       .op_out     (op_out_0_57),
       .pivot_out  (pivot_out_0_57),
       .r          (r_0_57)
     );

  // row 0, col 58

     reg start_in_0_58;
     wire start_out_0_58;

     reg swap_in_0_58;
     wire swap_out_0_58;

     reg [1:0] op_in_0_58;
     wire [1:0] op_out_0_58;

     wire r_0_58;

     wire data_in_0_58;
     wire data_out_0_58;

     reg pivot_in_0_58;
     wire pivot_out_0_58;

     assign data_in_0_58 = data_in[DAT_W-59];

     always @(posedge clk) begin
        op_in_0_58 <= op_out_0_57;
        pivot_in_0_58 <= pivot_out_0_57;
        start_in_0_58 <= start_out_0_57;
        swap_in_0_58 <= swap_out_0_57;
     end
  
     processor_AB AB_0_58 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_58),
       .start_in   (start_in_0_58),
       .swap_in    (swap_in_0_58),
       .op_in      (op_in_0_58),
       .pivot_in   (pivot_in_0_58),
       .start_out  (start_out_0_58),
       .swap_out   (swap_out_0_58),
       .data_out   (data_out_0_58),
       .op_out     (op_out_0_58),
       .pivot_out  (pivot_out_0_58),
       .r          (r_0_58)
     );

  // row 0, col 59

     reg start_in_0_59;
     wire start_out_0_59;

     reg swap_in_0_59;
     wire swap_out_0_59;

     reg [1:0] op_in_0_59;
     wire [1:0] op_out_0_59;

     wire r_0_59;

     wire data_in_0_59;
     wire data_out_0_59;

     reg pivot_in_0_59;
     wire pivot_out_0_59;

     assign data_in_0_59 = data_in[DAT_W-60];

     always @(posedge clk) begin
        op_in_0_59 <= op_out_0_58;
        pivot_in_0_59 <= pivot_out_0_58;
        start_in_0_59 <= start_out_0_58;
        swap_in_0_59 <= swap_out_0_58;
     end
  
     processor_AB AB_0_59 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_59),
       .start_in   (start_in_0_59),
       .swap_in    (swap_in_0_59),
       .op_in      (op_in_0_59),
       .pivot_in   (pivot_in_0_59),
       .start_out  (start_out_0_59),
       .swap_out   (swap_out_0_59),
       .data_out   (data_out_0_59),
       .op_out     (op_out_0_59),
       .pivot_out  (pivot_out_0_59),
       .r          (r_0_59)
     );

  // row 0, col 60

     reg start_in_0_60;
     wire start_out_0_60;

     reg swap_in_0_60;
     wire swap_out_0_60;

     reg [1:0] op_in_0_60;
     wire [1:0] op_out_0_60;

     wire r_0_60;

     wire data_in_0_60;
     wire data_out_0_60;

     reg pivot_in_0_60;
     wire pivot_out_0_60;

     assign data_in_0_60 = data_in[DAT_W-61];

     always @(posedge clk) begin
        op_in_0_60 <= op_out_0_59;
        pivot_in_0_60 <= pivot_out_0_59;
        start_in_0_60 <= start_out_0_59;
        swap_in_0_60 <= swap_out_0_59;
     end
  
     processor_AB AB_0_60 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_60),
       .start_in   (start_in_0_60),
       .swap_in    (swap_in_0_60),
       .op_in      (op_in_0_60),
       .pivot_in   (pivot_in_0_60),
       .start_out  (start_out_0_60),
       .swap_out   (swap_out_0_60),
       .data_out   (data_out_0_60),
       .op_out     (op_out_0_60),
       .pivot_out  (pivot_out_0_60),
       .r          (r_0_60)
     );

  // row 0, col 61

     reg start_in_0_61;
     wire start_out_0_61;

     reg swap_in_0_61;
     wire swap_out_0_61;

     reg [1:0] op_in_0_61;
     wire [1:0] op_out_0_61;

     wire r_0_61;

     wire data_in_0_61;
     wire data_out_0_61;

     reg pivot_in_0_61;
     wire pivot_out_0_61;

     assign data_in_0_61 = data_in[DAT_W-62];

     always @(posedge clk) begin
        op_in_0_61 <= op_out_0_60;
        pivot_in_0_61 <= pivot_out_0_60;
        start_in_0_61 <= start_out_0_60;
        swap_in_0_61 <= swap_out_0_60;
     end
  
     processor_AB AB_0_61 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_61),
       .start_in   (start_in_0_61),
       .swap_in    (swap_in_0_61),
       .op_in      (op_in_0_61),
       .pivot_in   (pivot_in_0_61),
       .start_out  (start_out_0_61),
       .swap_out   (swap_out_0_61),
       .data_out   (data_out_0_61),
       .op_out     (op_out_0_61),
       .pivot_out  (pivot_out_0_61),
       .r          (r_0_61)
     );

  // row 0, col 62

     reg start_in_0_62;
     wire start_out_0_62;

     reg swap_in_0_62;
     wire swap_out_0_62;

     reg [1:0] op_in_0_62;
     wire [1:0] op_out_0_62;

     wire r_0_62;

     wire data_in_0_62;
     wire data_out_0_62;

     reg pivot_in_0_62;
     wire pivot_out_0_62;

     assign data_in_0_62 = data_in[DAT_W-63];

     always @(posedge clk) begin
        op_in_0_62 <= op_out_0_61;
        pivot_in_0_62 <= pivot_out_0_61;
        start_in_0_62 <= start_out_0_61;
        swap_in_0_62 <= swap_out_0_61;
     end
  
     processor_AB AB_0_62 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_62),
       .start_in   (start_in_0_62),
       .swap_in    (swap_in_0_62),
       .op_in      (op_in_0_62),
       .pivot_in   (pivot_in_0_62),
       .start_out  (start_out_0_62),
       .swap_out   (swap_out_0_62),
       .data_out   (data_out_0_62),
       .op_out     (op_out_0_62),
       .pivot_out  (pivot_out_0_62),
       .r          (r_0_62)
     );

  // row 0, col 63

     reg start_in_0_63;
     wire start_out_0_63;

     reg swap_in_0_63;
     wire swap_out_0_63;

     reg [1:0] op_in_0_63;
     wire [1:0] op_out_0_63;

     wire r_0_63;

     wire data_in_0_63;
     wire data_out_0_63;

     reg pivot_in_0_63;
     wire pivot_out_0_63;

     assign data_in_0_63 = data_in[DAT_W-64];

     always @(posedge clk) begin
        op_in_0_63 <= op_out_0_62;
        pivot_in_0_63 <= pivot_out_0_62;
        start_in_0_63 <= start_out_0_62;
        swap_in_0_63 <= swap_out_0_62;
     end
  
     processor_AB AB_0_63 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_63),
       .start_in   (start_in_0_63),
       .swap_in    (swap_in_0_63),
       .op_in      (op_in_0_63),
       .pivot_in   (pivot_in_0_63),
       .start_out  (start_out_0_63),
       .swap_out   (swap_out_0_63),
       .data_out   (data_out_0_63),
       .op_out     (op_out_0_63),
       .pivot_out  (pivot_out_0_63),
       .r          (r_0_63)
     );

  // row 0, col 64

     reg start_in_0_64;
     wire start_out_0_64;

     reg swap_in_0_64;
     wire swap_out_0_64;

     reg [1:0] op_in_0_64;
     wire [1:0] op_out_0_64;

     wire r_0_64;

     wire data_in_0_64;
     wire data_out_0_64;

     reg pivot_in_0_64;
     wire pivot_out_0_64;

     assign data_in_0_64 = data_in[DAT_W-65];

     always @(posedge clk) begin
        op_in_0_64 <= op_out_0_63;
        pivot_in_0_64 <= pivot_out_0_63;
        start_in_0_64 <= start_out_0_63;
        swap_in_0_64 <= swap_out_0_63;
     end
  
     processor_AB AB_0_64 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_64),
       .start_in   (start_in_0_64),
       .swap_in    (swap_in_0_64),
       .op_in      (op_in_0_64),
       .pivot_in   (pivot_in_0_64),
       .start_out  (start_out_0_64),
       .swap_out   (swap_out_0_64),
       .data_out   (data_out_0_64),
       .op_out     (op_out_0_64),
       .pivot_out  (pivot_out_0_64),
       .r          (r_0_64)
     );

  // row 0, col 65

     reg start_in_0_65;
     wire start_out_0_65;

     reg swap_in_0_65;
     wire swap_out_0_65;

     reg [1:0] op_in_0_65;
     wire [1:0] op_out_0_65;

     wire r_0_65;

     wire data_in_0_65;
     wire data_out_0_65;

     reg pivot_in_0_65;
     wire pivot_out_0_65;

     assign data_in_0_65 = data_in[DAT_W-66];

     always @(posedge clk) begin
        op_in_0_65 <= op_out_0_64;
        pivot_in_0_65 <= pivot_out_0_64;
        start_in_0_65 <= start_out_0_64;
        swap_in_0_65 <= swap_out_0_64;
     end
  
     processor_AB AB_0_65 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_65),
       .start_in   (start_in_0_65),
       .swap_in    (swap_in_0_65),
       .op_in      (op_in_0_65),
       .pivot_in   (pivot_in_0_65),
       .start_out  (start_out_0_65),
       .swap_out   (swap_out_0_65),
       .data_out   (data_out_0_65),
       .op_out     (op_out_0_65),
       .pivot_out  (pivot_out_0_65),
       .r          (r_0_65)
     );

  // row 0, col 66

     reg start_in_0_66;
     wire start_out_0_66;

     reg swap_in_0_66;
     wire swap_out_0_66;

     reg [1:0] op_in_0_66;
     wire [1:0] op_out_0_66;

     wire r_0_66;

     wire data_in_0_66;
     wire data_out_0_66;

     reg pivot_in_0_66;
     wire pivot_out_0_66;

     assign data_in_0_66 = data_in[DAT_W-67];

     always @(posedge clk) begin
        op_in_0_66 <= op_out_0_65;
        pivot_in_0_66 <= pivot_out_0_65;
        start_in_0_66 <= start_out_0_65;
        swap_in_0_66 <= swap_out_0_65;
     end
  
     processor_AB AB_0_66 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_66),
       .start_in   (start_in_0_66),
       .swap_in    (swap_in_0_66),
       .op_in      (op_in_0_66),
       .pivot_in   (pivot_in_0_66),
       .start_out  (start_out_0_66),
       .swap_out   (swap_out_0_66),
       .data_out   (data_out_0_66),
       .op_out     (op_out_0_66),
       .pivot_out  (pivot_out_0_66),
       .r          (r_0_66)
     );

  // row 0, col 67

     reg start_in_0_67;
     wire start_out_0_67;

     reg swap_in_0_67;
     wire swap_out_0_67;

     reg [1:0] op_in_0_67;
     wire [1:0] op_out_0_67;

     wire r_0_67;

     wire data_in_0_67;
     wire data_out_0_67;

     reg pivot_in_0_67;
     wire pivot_out_0_67;

     assign data_in_0_67 = data_in[DAT_W-68];

     always @(posedge clk) begin
        op_in_0_67 <= op_out_0_66;
        pivot_in_0_67 <= pivot_out_0_66;
        start_in_0_67 <= start_out_0_66;
        swap_in_0_67 <= swap_out_0_66;
     end
  
     processor_AB AB_0_67 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_67),
       .start_in   (start_in_0_67),
       .swap_in    (swap_in_0_67),
       .op_in      (op_in_0_67),
       .pivot_in   (pivot_in_0_67),
       .start_out  (start_out_0_67),
       .swap_out   (swap_out_0_67),
       .data_out   (data_out_0_67),
       .op_out     (op_out_0_67),
       .pivot_out  (pivot_out_0_67),
       .r          (r_0_67)
     );

  // row 0, col 68

     reg start_in_0_68;
     wire start_out_0_68;

     reg swap_in_0_68;
     wire swap_out_0_68;

     reg [1:0] op_in_0_68;
     wire [1:0] op_out_0_68;

     wire r_0_68;

     wire data_in_0_68;
     wire data_out_0_68;

     reg pivot_in_0_68;
     wire pivot_out_0_68;

     assign data_in_0_68 = data_in[DAT_W-69];

     always @(posedge clk) begin
        op_in_0_68 <= op_out_0_67;
        pivot_in_0_68 <= pivot_out_0_67;
        start_in_0_68 <= start_out_0_67;
        swap_in_0_68 <= swap_out_0_67;
     end
  
     processor_AB AB_0_68 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_68),
       .start_in   (start_in_0_68),
       .swap_in    (swap_in_0_68),
       .op_in      (op_in_0_68),
       .pivot_in   (pivot_in_0_68),
       .start_out  (start_out_0_68),
       .swap_out   (swap_out_0_68),
       .data_out   (data_out_0_68),
       .op_out     (op_out_0_68),
       .pivot_out  (pivot_out_0_68),
       .r          (r_0_68)
     );

  // row 0, col 69

     reg start_in_0_69;
     wire start_out_0_69;

     reg swap_in_0_69;
     wire swap_out_0_69;

     reg [1:0] op_in_0_69;
     wire [1:0] op_out_0_69;

     wire r_0_69;

     wire data_in_0_69;
     wire data_out_0_69;

     reg pivot_in_0_69;
     wire pivot_out_0_69;

     assign data_in_0_69 = data_in[DAT_W-70];

     always @(posedge clk) begin
        op_in_0_69 <= op_out_0_68;
        pivot_in_0_69 <= pivot_out_0_68;
        start_in_0_69 <= start_out_0_68;
        swap_in_0_69 <= swap_out_0_68;
     end
  
     processor_AB AB_0_69 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_69),
       .start_in   (start_in_0_69),
       .swap_in    (swap_in_0_69),
       .op_in      (op_in_0_69),
       .pivot_in   (pivot_in_0_69),
       .start_out  (start_out_0_69),
       .swap_out   (swap_out_0_69),
       .data_out   (data_out_0_69),
       .op_out     (op_out_0_69),
       .pivot_out  (pivot_out_0_69),
       .r          (r_0_69)
     );

  // row 0, col 70

     reg start_in_0_70;
     wire start_out_0_70;

     reg swap_in_0_70;
     wire swap_out_0_70;

     reg [1:0] op_in_0_70;
     wire [1:0] op_out_0_70;

     wire r_0_70;

     wire data_in_0_70;
     wire data_out_0_70;

     reg pivot_in_0_70;
     wire pivot_out_0_70;

     assign data_in_0_70 = data_in[DAT_W-71];

     always @(posedge clk) begin
        op_in_0_70 <= op_out_0_69;
        pivot_in_0_70 <= pivot_out_0_69;
        start_in_0_70 <= start_out_0_69;
        swap_in_0_70 <= swap_out_0_69;
     end
  
     processor_AB AB_0_70 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_70),
       .start_in   (start_in_0_70),
       .swap_in    (swap_in_0_70),
       .op_in      (op_in_0_70),
       .pivot_in   (pivot_in_0_70),
       .start_out  (start_out_0_70),
       .swap_out   (swap_out_0_70),
       .data_out   (data_out_0_70),
       .op_out     (op_out_0_70),
       .pivot_out  (pivot_out_0_70),
       .r          (r_0_70)
     );

  // row 0, col 71

     reg start_in_0_71;
     wire start_out_0_71;

     reg swap_in_0_71;
     wire swap_out_0_71;

     reg [1:0] op_in_0_71;
     wire [1:0] op_out_0_71;

     wire r_0_71;

     wire data_in_0_71;
     wire data_out_0_71;

     reg pivot_in_0_71;
     wire pivot_out_0_71;

     assign data_in_0_71 = data_in[DAT_W-72];

     always @(posedge clk) begin
        op_in_0_71 <= op_out_0_70;
        pivot_in_0_71 <= pivot_out_0_70;
        start_in_0_71 <= start_out_0_70;
        swap_in_0_71 <= swap_out_0_70;
     end
  
     processor_AB AB_0_71 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_71),
       .start_in   (start_in_0_71),
       .swap_in    (swap_in_0_71),
       .op_in      (op_in_0_71),
       .pivot_in   (pivot_in_0_71),
       .start_out  (start_out_0_71),
       .swap_out   (swap_out_0_71),
       .data_out   (data_out_0_71),
       .op_out     (op_out_0_71),
       .pivot_out  (pivot_out_0_71),
       .r          (r_0_71)
     );

  // row 0, col 72

     reg start_in_0_72;
     wire start_out_0_72;

     reg swap_in_0_72;
     wire swap_out_0_72;

     reg [1:0] op_in_0_72;
     wire [1:0] op_out_0_72;

     wire r_0_72;

     wire data_in_0_72;
     wire data_out_0_72;

     reg pivot_in_0_72;
     wire pivot_out_0_72;

     assign data_in_0_72 = data_in[DAT_W-73];

     always @(posedge clk) begin
        op_in_0_72 <= op_out_0_71;
        pivot_in_0_72 <= pivot_out_0_71;
        start_in_0_72 <= start_out_0_71;
        swap_in_0_72 <= swap_out_0_71;
     end
  
     processor_AB AB_0_72 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_72),
       .start_in   (start_in_0_72),
       .swap_in    (swap_in_0_72),
       .op_in      (op_in_0_72),
       .pivot_in   (pivot_in_0_72),
       .start_out  (start_out_0_72),
       .swap_out   (swap_out_0_72),
       .data_out   (data_out_0_72),
       .op_out     (op_out_0_72),
       .pivot_out  (pivot_out_0_72),
       .r          (r_0_72)
     );

  // row 0, col 73

     reg start_in_0_73;
     wire start_out_0_73;

     reg swap_in_0_73;
     wire swap_out_0_73;

     reg [1:0] op_in_0_73;
     wire [1:0] op_out_0_73;

     wire r_0_73;

     wire data_in_0_73;
     wire data_out_0_73;

     reg pivot_in_0_73;
     wire pivot_out_0_73;

     assign data_in_0_73 = data_in[DAT_W-74];

     always @(posedge clk) begin
        op_in_0_73 <= op_out_0_72;
        pivot_in_0_73 <= pivot_out_0_72;
        start_in_0_73 <= start_out_0_72;
        swap_in_0_73 <= swap_out_0_72;
     end
  
     processor_AB AB_0_73 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_73),
       .start_in   (start_in_0_73),
       .swap_in    (swap_in_0_73),
       .op_in      (op_in_0_73),
       .pivot_in   (pivot_in_0_73),
       .start_out  (start_out_0_73),
       .swap_out   (swap_out_0_73),
       .data_out   (data_out_0_73),
       .op_out     (op_out_0_73),
       .pivot_out  (pivot_out_0_73),
       .r          (r_0_73)
     );

  // row 0, col 74

     reg start_in_0_74;
     wire start_out_0_74;

     reg swap_in_0_74;
     wire swap_out_0_74;

     reg [1:0] op_in_0_74;
     wire [1:0] op_out_0_74;

     wire r_0_74;

     wire data_in_0_74;
     wire data_out_0_74;

     reg pivot_in_0_74;
     wire pivot_out_0_74;

     assign data_in_0_74 = data_in[DAT_W-75];

     always @(posedge clk) begin
        op_in_0_74 <= op_out_0_73;
        pivot_in_0_74 <= pivot_out_0_73;
        start_in_0_74 <= start_out_0_73;
        swap_in_0_74 <= swap_out_0_73;
     end
  
     processor_AB AB_0_74 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_74),
       .start_in   (start_in_0_74),
       .swap_in    (swap_in_0_74),
       .op_in      (op_in_0_74),
       .pivot_in   (pivot_in_0_74),
       .start_out  (start_out_0_74),
       .swap_out   (swap_out_0_74),
       .data_out   (data_out_0_74),
       .op_out     (op_out_0_74),
       .pivot_out  (pivot_out_0_74),
       .r          (r_0_74)
     );

  // row 0, col 75

     reg start_in_0_75;
     wire start_out_0_75;

     reg swap_in_0_75;
     wire swap_out_0_75;

     reg [1:0] op_in_0_75;
     wire [1:0] op_out_0_75;

     wire r_0_75;

     wire data_in_0_75;
     wire data_out_0_75;

     reg pivot_in_0_75;
     wire pivot_out_0_75;

     assign data_in_0_75 = data_in[DAT_W-76];

     always @(posedge clk) begin
        op_in_0_75 <= op_out_0_74;
        pivot_in_0_75 <= pivot_out_0_74;
        start_in_0_75 <= start_out_0_74;
        swap_in_0_75 <= swap_out_0_74;
     end
  
     processor_AB AB_0_75 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_75),
       .start_in   (start_in_0_75),
       .swap_in    (swap_in_0_75),
       .op_in      (op_in_0_75),
       .pivot_in   (pivot_in_0_75),
       .start_out  (start_out_0_75),
       .swap_out   (swap_out_0_75),
       .data_out   (data_out_0_75),
       .op_out     (op_out_0_75),
       .pivot_out  (pivot_out_0_75),
       .r          (r_0_75)
     );

  // row 0, col 76

     reg start_in_0_76;
     wire start_out_0_76;

     reg swap_in_0_76;
     wire swap_out_0_76;

     reg [1:0] op_in_0_76;
     wire [1:0] op_out_0_76;

     wire r_0_76;

     wire data_in_0_76;
     wire data_out_0_76;

     reg pivot_in_0_76;
     wire pivot_out_0_76;

     assign data_in_0_76 = data_in[DAT_W-77];

     always @(posedge clk) begin
        op_in_0_76 <= op_out_0_75;
        pivot_in_0_76 <= pivot_out_0_75;
        start_in_0_76 <= start_out_0_75;
        swap_in_0_76 <= swap_out_0_75;
     end
  
     processor_AB AB_0_76 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_76),
       .start_in   (start_in_0_76),
       .swap_in    (swap_in_0_76),
       .op_in      (op_in_0_76),
       .pivot_in   (pivot_in_0_76),
       .start_out  (start_out_0_76),
       .swap_out   (swap_out_0_76),
       .data_out   (data_out_0_76),
       .op_out     (op_out_0_76),
       .pivot_out  (pivot_out_0_76),
       .r          (r_0_76)
     );

  // row 0, col 77

     reg start_in_0_77;
     wire start_out_0_77;

     reg swap_in_0_77;
     wire swap_out_0_77;

     reg [1:0] op_in_0_77;
     wire [1:0] op_out_0_77;

     wire r_0_77;

     wire data_in_0_77;
     wire data_out_0_77;

     reg pivot_in_0_77;
     wire pivot_out_0_77;

     assign data_in_0_77 = data_in[DAT_W-78];

     always @(posedge clk) begin
        op_in_0_77 <= op_out_0_76;
        pivot_in_0_77 <= pivot_out_0_76;
        start_in_0_77 <= start_out_0_76;
        swap_in_0_77 <= swap_out_0_76;
     end
  
     processor_AB AB_0_77 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_77),
       .start_in   (start_in_0_77),
       .swap_in    (swap_in_0_77),
       .op_in      (op_in_0_77),
       .pivot_in   (pivot_in_0_77),
       .start_out  (start_out_0_77),
       .swap_out   (swap_out_0_77),
       .data_out   (data_out_0_77),
       .op_out     (op_out_0_77),
       .pivot_out  (pivot_out_0_77),
       .r          (r_0_77)
     );

  // row 0, col 78

     reg start_in_0_78;
     wire start_out_0_78;

     reg swap_in_0_78;
     wire swap_out_0_78;

     reg [1:0] op_in_0_78;
     wire [1:0] op_out_0_78;

     wire r_0_78;

     wire data_in_0_78;
     wire data_out_0_78;

     reg pivot_in_0_78;
     wire pivot_out_0_78;

     assign data_in_0_78 = data_in[DAT_W-79];

     always @(posedge clk) begin
        op_in_0_78 <= op_out_0_77;
        pivot_in_0_78 <= pivot_out_0_77;
        start_in_0_78 <= start_out_0_77;
        swap_in_0_78 <= swap_out_0_77;
     end
  
     processor_AB AB_0_78 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_78),
       .start_in   (start_in_0_78),
       .swap_in    (swap_in_0_78),
       .op_in      (op_in_0_78),
       .pivot_in   (pivot_in_0_78),
       .start_out  (start_out_0_78),
       .swap_out   (swap_out_0_78),
       .data_out   (data_out_0_78),
       .op_out     (op_out_0_78),
       .pivot_out  (pivot_out_0_78),
       .r          (r_0_78)
     );

  // row 0, col 79

     reg start_in_0_79;
     wire start_out_0_79;

     reg swap_in_0_79;
     wire swap_out_0_79;

     reg [1:0] op_in_0_79;
     wire [1:0] op_out_0_79;

     wire r_0_79;

     wire data_in_0_79;
     wire data_out_0_79;

     reg pivot_in_0_79;
     wire pivot_out_0_79;

     assign data_in_0_79 = data_in[DAT_W-80];

     always @(posedge clk) begin
        op_in_0_79 <= op_out_0_78;
        pivot_in_0_79 <= pivot_out_0_78;
        start_in_0_79 <= start_out_0_78;
        swap_in_0_79 <= swap_out_0_78;
     end
  
     processor_AB AB_0_79 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_79),
       .start_in   (start_in_0_79),
       .swap_in    (swap_in_0_79),
       .op_in      (op_in_0_79),
       .pivot_in   (pivot_in_0_79),
       .start_out  (start_out_0_79),
       .swap_out   (swap_out_0_79),
       .data_out   (data_out_0_79),
       .op_out     (op_out_0_79),
       .pivot_out  (pivot_out_0_79),
       .r          (r_0_79)
     );

  // row 0, col 80

     reg start_in_0_80;
     wire start_out_0_80;

     reg swap_in_0_80;
     wire swap_out_0_80;

     reg [1:0] op_in_0_80;
     wire [1:0] op_out_0_80;

     wire r_0_80;

     wire data_in_0_80;
     wire data_out_0_80;

     reg pivot_in_0_80;
     wire pivot_out_0_80;

     assign data_in_0_80 = data_in[DAT_W-81];

     always @(posedge clk) begin
        op_in_0_80 <= op_out_0_79;
        pivot_in_0_80 <= pivot_out_0_79;
        start_in_0_80 <= start_out_0_79;
        swap_in_0_80 <= swap_out_0_79;
     end
  
     processor_AB AB_0_80 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_80),
       .start_in   (start_in_0_80),
       .swap_in    (swap_in_0_80),
       .op_in      (op_in_0_80),
       .pivot_in   (pivot_in_0_80),
       .start_out  (start_out_0_80),
       .swap_out   (swap_out_0_80),
       .data_out   (data_out_0_80),
       .op_out     (op_out_0_80),
       .pivot_out  (pivot_out_0_80),
       .r          (r_0_80)
     );

  // row 0, col 81

     reg start_in_0_81;
     wire start_out_0_81;

     reg swap_in_0_81;
     wire swap_out_0_81;

     reg [1:0] op_in_0_81;
     wire [1:0] op_out_0_81;

     wire r_0_81;

     wire data_in_0_81;
     wire data_out_0_81;

     reg pivot_in_0_81;
     wire pivot_out_0_81;

     assign data_in_0_81 = data_in[DAT_W-82];

     always @(posedge clk) begin
        op_in_0_81 <= op_out_0_80;
        pivot_in_0_81 <= pivot_out_0_80;
        start_in_0_81 <= start_out_0_80;
        swap_in_0_81 <= swap_out_0_80;
     end
  
     processor_AB AB_0_81 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_81),
       .start_in   (start_in_0_81),
       .swap_in    (swap_in_0_81),
       .op_in      (op_in_0_81),
       .pivot_in   (pivot_in_0_81),
       .start_out  (start_out_0_81),
       .swap_out   (swap_out_0_81),
       .data_out   (data_out_0_81),
       .op_out     (op_out_0_81),
       .pivot_out  (pivot_out_0_81),
       .r          (r_0_81)
     );

  // row 0, col 82

     reg start_in_0_82;
     wire start_out_0_82;

     reg swap_in_0_82;
     wire swap_out_0_82;

     reg [1:0] op_in_0_82;
     wire [1:0] op_out_0_82;

     wire r_0_82;

     wire data_in_0_82;
     wire data_out_0_82;

     reg pivot_in_0_82;
     wire pivot_out_0_82;

     assign data_in_0_82 = data_in[DAT_W-83];

     always @(posedge clk) begin
        op_in_0_82 <= op_out_0_81;
        pivot_in_0_82 <= pivot_out_0_81;
        start_in_0_82 <= start_out_0_81;
        swap_in_0_82 <= swap_out_0_81;
     end
  
     processor_AB AB_0_82 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_82),
       .start_in   (start_in_0_82),
       .swap_in    (swap_in_0_82),
       .op_in      (op_in_0_82),
       .pivot_in   (pivot_in_0_82),
       .start_out  (start_out_0_82),
       .swap_out   (swap_out_0_82),
       .data_out   (data_out_0_82),
       .op_out     (op_out_0_82),
       .pivot_out  (pivot_out_0_82),
       .r          (r_0_82)
     );

  // row 0, col 83

     reg start_in_0_83;
     wire start_out_0_83;

     reg swap_in_0_83;
     wire swap_out_0_83;

     reg [1:0] op_in_0_83;
     wire [1:0] op_out_0_83;

     wire r_0_83;

     wire data_in_0_83;
     wire data_out_0_83;

     reg pivot_in_0_83;
     wire pivot_out_0_83;

     assign data_in_0_83 = data_in[DAT_W-84];

     always @(posedge clk) begin
        op_in_0_83 <= op_out_0_82;
        pivot_in_0_83 <= pivot_out_0_82;
        start_in_0_83 <= start_out_0_82;
        swap_in_0_83 <= swap_out_0_82;
     end
  
     processor_AB AB_0_83 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_83),
       .start_in   (start_in_0_83),
       .swap_in    (swap_in_0_83),
       .op_in      (op_in_0_83),
       .pivot_in   (pivot_in_0_83),
       .start_out  (start_out_0_83),
       .swap_out   (swap_out_0_83),
       .data_out   (data_out_0_83),
       .op_out     (op_out_0_83),
       .pivot_out  (pivot_out_0_83),
       .r          (r_0_83)
     );

  // row 0, col 84

     reg start_in_0_84;
     wire start_out_0_84;

     reg swap_in_0_84;
     wire swap_out_0_84;

     reg [1:0] op_in_0_84;
     wire [1:0] op_out_0_84;

     wire r_0_84;

     wire data_in_0_84;
     wire data_out_0_84;

     reg pivot_in_0_84;
     wire pivot_out_0_84;

     assign data_in_0_84 = data_in[DAT_W-85];

     always @(posedge clk) begin
        op_in_0_84 <= op_out_0_83;
        pivot_in_0_84 <= pivot_out_0_83;
        start_in_0_84 <= start_out_0_83;
        swap_in_0_84 <= swap_out_0_83;
     end
  
     processor_AB AB_0_84 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_84),
       .start_in   (start_in_0_84),
       .swap_in    (swap_in_0_84),
       .op_in      (op_in_0_84),
       .pivot_in   (pivot_in_0_84),
       .start_out  (start_out_0_84),
       .swap_out   (swap_out_0_84),
       .data_out   (data_out_0_84),
       .op_out     (op_out_0_84),
       .pivot_out  (pivot_out_0_84),
       .r          (r_0_84)
     );

  // row 0, col 85

     reg start_in_0_85;
     wire start_out_0_85;

     reg swap_in_0_85;
     wire swap_out_0_85;

     reg [1:0] op_in_0_85;
     wire [1:0] op_out_0_85;

     wire r_0_85;

     wire data_in_0_85;
     wire data_out_0_85;

     reg pivot_in_0_85;
     wire pivot_out_0_85;

     assign data_in_0_85 = data_in[DAT_W-86];

     always @(posedge clk) begin
        op_in_0_85 <= op_out_0_84;
        pivot_in_0_85 <= pivot_out_0_84;
        start_in_0_85 <= start_out_0_84;
        swap_in_0_85 <= swap_out_0_84;
     end
  
     processor_AB AB_0_85 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_85),
       .start_in   (start_in_0_85),
       .swap_in    (swap_in_0_85),
       .op_in      (op_in_0_85),
       .pivot_in   (pivot_in_0_85),
       .start_out  (start_out_0_85),
       .swap_out   (swap_out_0_85),
       .data_out   (data_out_0_85),
       .op_out     (op_out_0_85),
       .pivot_out  (pivot_out_0_85),
       .r          (r_0_85)
     );

  // row 0, col 86

     reg start_in_0_86;
     wire start_out_0_86;

     reg swap_in_0_86;
     wire swap_out_0_86;

     reg [1:0] op_in_0_86;
     wire [1:0] op_out_0_86;

     wire r_0_86;

     wire data_in_0_86;
     wire data_out_0_86;

     reg pivot_in_0_86;
     wire pivot_out_0_86;

     assign data_in_0_86 = data_in[DAT_W-87];

     always @(posedge clk) begin
        op_in_0_86 <= op_out_0_85;
        pivot_in_0_86 <= pivot_out_0_85;
        start_in_0_86 <= start_out_0_85;
        swap_in_0_86 <= swap_out_0_85;
     end
  
     processor_AB AB_0_86 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_86),
       .start_in   (start_in_0_86),
       .swap_in    (swap_in_0_86),
       .op_in      (op_in_0_86),
       .pivot_in   (pivot_in_0_86),
       .start_out  (start_out_0_86),
       .swap_out   (swap_out_0_86),
       .data_out   (data_out_0_86),
       .op_out     (op_out_0_86),
       .pivot_out  (pivot_out_0_86),
       .r          (r_0_86)
     );

  // row 0, col 87

     reg start_in_0_87;
     wire start_out_0_87;

     reg swap_in_0_87;
     wire swap_out_0_87;

     reg [1:0] op_in_0_87;
     wire [1:0] op_out_0_87;

     wire r_0_87;

     wire data_in_0_87;
     wire data_out_0_87;

     reg pivot_in_0_87;
     wire pivot_out_0_87;

     assign data_in_0_87 = data_in[DAT_W-88];

     always @(posedge clk) begin
        op_in_0_87 <= op_out_0_86;
        pivot_in_0_87 <= pivot_out_0_86;
        start_in_0_87 <= start_out_0_86;
        swap_in_0_87 <= swap_out_0_86;
     end
  
     processor_AB AB_0_87 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_87),
       .start_in   (start_in_0_87),
       .swap_in    (swap_in_0_87),
       .op_in      (op_in_0_87),
       .pivot_in   (pivot_in_0_87),
       .start_out  (start_out_0_87),
       .swap_out   (swap_out_0_87),
       .data_out   (data_out_0_87),
       .op_out     (op_out_0_87),
       .pivot_out  (pivot_out_0_87),
       .r          (r_0_87)
     );

  // row 0, col 88

     reg start_in_0_88;
     wire start_out_0_88;

     reg swap_in_0_88;
     wire swap_out_0_88;

     reg [1:0] op_in_0_88;
     wire [1:0] op_out_0_88;

     wire r_0_88;

     wire data_in_0_88;
     wire data_out_0_88;

     reg pivot_in_0_88;
     wire pivot_out_0_88;

     assign data_in_0_88 = data_in[DAT_W-89];

     always @(posedge clk) begin
        op_in_0_88 <= op_out_0_87;
        pivot_in_0_88 <= pivot_out_0_87;
        start_in_0_88 <= start_out_0_87;
        swap_in_0_88 <= swap_out_0_87;
     end
  
     processor_AB AB_0_88 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_88),
       .start_in   (start_in_0_88),
       .swap_in    (swap_in_0_88),
       .op_in      (op_in_0_88),
       .pivot_in   (pivot_in_0_88),
       .start_out  (start_out_0_88),
       .swap_out   (swap_out_0_88),
       .data_out   (data_out_0_88),
       .op_out     (op_out_0_88),
       .pivot_out  (pivot_out_0_88),
       .r          (r_0_88)
     );

  // row 0, col 89

     reg start_in_0_89;
     wire start_out_0_89;

     reg swap_in_0_89;
     wire swap_out_0_89;

     reg [1:0] op_in_0_89;
     wire [1:0] op_out_0_89;

     wire r_0_89;

     wire data_in_0_89;
     wire data_out_0_89;

     reg pivot_in_0_89;
     wire pivot_out_0_89;

     assign data_in_0_89 = data_in[DAT_W-90];

     always @(posedge clk) begin
        op_in_0_89 <= op_out_0_88;
        pivot_in_0_89 <= pivot_out_0_88;
        start_in_0_89 <= start_out_0_88;
        swap_in_0_89 <= swap_out_0_88;
     end
  
     processor_AB AB_0_89 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_89),
       .start_in   (start_in_0_89),
       .swap_in    (swap_in_0_89),
       .op_in      (op_in_0_89),
       .pivot_in   (pivot_in_0_89),
       .start_out  (start_out_0_89),
       .swap_out   (swap_out_0_89),
       .data_out   (data_out_0_89),
       .op_out     (op_out_0_89),
       .pivot_out  (pivot_out_0_89),
       .r          (r_0_89)
     );

  // row 0, col 90

     reg start_in_0_90;
     wire start_out_0_90;

     reg swap_in_0_90;
     wire swap_out_0_90;

     reg [1:0] op_in_0_90;
     wire [1:0] op_out_0_90;

     wire r_0_90;

     wire data_in_0_90;
     wire data_out_0_90;

     reg pivot_in_0_90;
     wire pivot_out_0_90;

     assign data_in_0_90 = data_in[DAT_W-91];

     always @(posedge clk) begin
        op_in_0_90 <= op_out_0_89;
        pivot_in_0_90 <= pivot_out_0_89;
        start_in_0_90 <= start_out_0_89;
        swap_in_0_90 <= swap_out_0_89;
     end
  
     processor_AB AB_0_90 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_90),
       .start_in   (start_in_0_90),
       .swap_in    (swap_in_0_90),
       .op_in      (op_in_0_90),
       .pivot_in   (pivot_in_0_90),
       .start_out  (start_out_0_90),
       .swap_out   (swap_out_0_90),
       .data_out   (data_out_0_90),
       .op_out     (op_out_0_90),
       .pivot_out  (pivot_out_0_90),
       .r          (r_0_90)
     );

  // row 0, col 91

     reg start_in_0_91;
     wire start_out_0_91;

     reg swap_in_0_91;
     wire swap_out_0_91;

     reg [1:0] op_in_0_91;
     wire [1:0] op_out_0_91;

     wire r_0_91;

     wire data_in_0_91;
     wire data_out_0_91;

     reg pivot_in_0_91;
     wire pivot_out_0_91;

     assign data_in_0_91 = data_in[DAT_W-92];

     always @(posedge clk) begin
        op_in_0_91 <= op_out_0_90;
        pivot_in_0_91 <= pivot_out_0_90;
        start_in_0_91 <= start_out_0_90;
        swap_in_0_91 <= swap_out_0_90;
     end
  
     processor_AB AB_0_91 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_91),
       .start_in   (start_in_0_91),
       .swap_in    (swap_in_0_91),
       .op_in      (op_in_0_91),
       .pivot_in   (pivot_in_0_91),
       .start_out  (start_out_0_91),
       .swap_out   (swap_out_0_91),
       .data_out   (data_out_0_91),
       .op_out     (op_out_0_91),
       .pivot_out  (pivot_out_0_91),
       .r          (r_0_91)
     );

  // row 0, col 92

     reg start_in_0_92;
     wire start_out_0_92;

     reg swap_in_0_92;
     wire swap_out_0_92;

     reg [1:0] op_in_0_92;
     wire [1:0] op_out_0_92;

     wire r_0_92;

     wire data_in_0_92;
     wire data_out_0_92;

     reg pivot_in_0_92;
     wire pivot_out_0_92;

     assign data_in_0_92 = data_in[DAT_W-93];

     always @(posedge clk) begin
        op_in_0_92 <= op_out_0_91;
        pivot_in_0_92 <= pivot_out_0_91;
        start_in_0_92 <= start_out_0_91;
        swap_in_0_92 <= swap_out_0_91;
     end
  
     processor_AB AB_0_92 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_92),
       .start_in   (start_in_0_92),
       .swap_in    (swap_in_0_92),
       .op_in      (op_in_0_92),
       .pivot_in   (pivot_in_0_92),
       .start_out  (start_out_0_92),
       .swap_out   (swap_out_0_92),
       .data_out   (data_out_0_92),
       .op_out     (op_out_0_92),
       .pivot_out  (pivot_out_0_92),
       .r          (r_0_92)
     );

  // row 0, col 93

     reg start_in_0_93;
     wire start_out_0_93;

     reg swap_in_0_93;
     wire swap_out_0_93;

     reg [1:0] op_in_0_93;
     wire [1:0] op_out_0_93;

     wire r_0_93;

     wire data_in_0_93;
     wire data_out_0_93;

     reg pivot_in_0_93;
     wire pivot_out_0_93;

     assign data_in_0_93 = data_in[DAT_W-94];

     always @(posedge clk) begin
        op_in_0_93 <= op_out_0_92;
        pivot_in_0_93 <= pivot_out_0_92;
        start_in_0_93 <= start_out_0_92;
        swap_in_0_93 <= swap_out_0_92;
     end
  
     processor_AB AB_0_93 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_93),
       .start_in   (start_in_0_93),
       .swap_in    (swap_in_0_93),
       .op_in      (op_in_0_93),
       .pivot_in   (pivot_in_0_93),
       .start_out  (start_out_0_93),
       .swap_out   (swap_out_0_93),
       .data_out   (data_out_0_93),
       .op_out     (op_out_0_93),
       .pivot_out  (pivot_out_0_93),
       .r          (r_0_93)
     );

  // row 0, col 94

     reg start_in_0_94;
     wire start_out_0_94;

     reg swap_in_0_94;
     wire swap_out_0_94;

     reg [1:0] op_in_0_94;
     wire [1:0] op_out_0_94;

     wire r_0_94;

     wire data_in_0_94;
     wire data_out_0_94;

     reg pivot_in_0_94;
     wire pivot_out_0_94;

     assign data_in_0_94 = data_in[DAT_W-95];

     always @(posedge clk) begin
        op_in_0_94 <= op_out_0_93;
        pivot_in_0_94 <= pivot_out_0_93;
        start_in_0_94 <= start_out_0_93;
        swap_in_0_94 <= swap_out_0_93;
     end
  
     processor_AB AB_0_94 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_94),
       .start_in   (start_in_0_94),
       .swap_in    (swap_in_0_94),
       .op_in      (op_in_0_94),
       .pivot_in   (pivot_in_0_94),
       .start_out  (start_out_0_94),
       .swap_out   (swap_out_0_94),
       .data_out   (data_out_0_94),
       .op_out     (op_out_0_94),
       .pivot_out  (pivot_out_0_94),
       .r          (r_0_94)
     );

  // row 0, col 95

     reg start_in_0_95;
     wire start_out_0_95;

     reg swap_in_0_95;
     wire swap_out_0_95;

     reg [1:0] op_in_0_95;
     wire [1:0] op_out_0_95;

     wire r_0_95;

     wire data_in_0_95;
     wire data_out_0_95;

     reg pivot_in_0_95;
     wire pivot_out_0_95;

     assign data_in_0_95 = data_in[DAT_W-96];

     always @(posedge clk) begin
        op_in_0_95 <= op_out_0_94;
        pivot_in_0_95 <= pivot_out_0_94;
        start_in_0_95 <= start_out_0_94;
        swap_in_0_95 <= swap_out_0_94;
     end
  
     processor_AB AB_0_95 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_95),
       .start_in   (start_in_0_95),
       .swap_in    (swap_in_0_95),
       .op_in      (op_in_0_95),
       .pivot_in   (pivot_in_0_95),
       .start_out  (start_out_0_95),
       .swap_out   (swap_out_0_95),
       .data_out   (data_out_0_95),
       .op_out     (op_out_0_95),
       .pivot_out  (pivot_out_0_95),
       .r          (r_0_95)
     );

  // row 0, col 96

     reg start_in_0_96;
     wire start_out_0_96;

     reg swap_in_0_96;
     wire swap_out_0_96;

     reg [1:0] op_in_0_96;
     wire [1:0] op_out_0_96;

     wire r_0_96;

     wire data_in_0_96;
     wire data_out_0_96;

     reg pivot_in_0_96;
     wire pivot_out_0_96;

     assign data_in_0_96 = data_in[DAT_W-97];

     always @(posedge clk) begin
        op_in_0_96 <= op_out_0_95;
        pivot_in_0_96 <= pivot_out_0_95;
        start_in_0_96 <= start_out_0_95;
        swap_in_0_96 <= swap_out_0_95;
     end
  
     processor_AB AB_0_96 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_96),
       .start_in   (start_in_0_96),
       .swap_in    (swap_in_0_96),
       .op_in      (op_in_0_96),
       .pivot_in   (pivot_in_0_96),
       .start_out  (start_out_0_96),
       .swap_out   (swap_out_0_96),
       .data_out   (data_out_0_96),
       .op_out     (op_out_0_96),
       .pivot_out  (pivot_out_0_96),
       .r          (r_0_96)
     );

  // row 0, col 97

     reg start_in_0_97;
     wire start_out_0_97;

     reg swap_in_0_97;
     wire swap_out_0_97;

     reg [1:0] op_in_0_97;
     wire [1:0] op_out_0_97;

     wire r_0_97;

     wire data_in_0_97;
     wire data_out_0_97;

     reg pivot_in_0_97;
     wire pivot_out_0_97;

     assign data_in_0_97 = data_in[DAT_W-98];

     always @(posedge clk) begin
        op_in_0_97 <= op_out_0_96;
        pivot_in_0_97 <= pivot_out_0_96;
        start_in_0_97 <= start_out_0_96;
        swap_in_0_97 <= swap_out_0_96;
     end
  
     processor_AB AB_0_97 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_97),
       .start_in   (start_in_0_97),
       .swap_in    (swap_in_0_97),
       .op_in      (op_in_0_97),
       .pivot_in   (pivot_in_0_97),
       .start_out  (start_out_0_97),
       .swap_out   (swap_out_0_97),
       .data_out   (data_out_0_97),
       .op_out     (op_out_0_97),
       .pivot_out  (pivot_out_0_97),
       .r          (r_0_97)
     );

  // row 0, col 98

     reg start_in_0_98;
     wire start_out_0_98;

     reg swap_in_0_98;
     wire swap_out_0_98;

     reg [1:0] op_in_0_98;
     wire [1:0] op_out_0_98;

     wire r_0_98;

     wire data_in_0_98;
     wire data_out_0_98;

     reg pivot_in_0_98;
     wire pivot_out_0_98;

     assign data_in_0_98 = data_in[DAT_W-99];

     always @(posedge clk) begin
        op_in_0_98 <= op_out_0_97;
        pivot_in_0_98 <= pivot_out_0_97;
        start_in_0_98 <= start_out_0_97;
        swap_in_0_98 <= swap_out_0_97;
     end
  
     processor_AB AB_0_98 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_98),
       .start_in   (start_in_0_98),
       .swap_in    (swap_in_0_98),
       .op_in      (op_in_0_98),
       .pivot_in   (pivot_in_0_98),
       .start_out  (start_out_0_98),
       .swap_out   (swap_out_0_98),
       .data_out   (data_out_0_98),
       .op_out     (op_out_0_98),
       .pivot_out  (pivot_out_0_98),
       .r          (r_0_98)
     );

  // row 0, col 99

     reg start_in_0_99;
     wire start_out_0_99;

     reg swap_in_0_99;
     wire swap_out_0_99;

     reg [1:0] op_in_0_99;
     wire [1:0] op_out_0_99;

     wire r_0_99;

     wire data_in_0_99;
     wire data_out_0_99;

     reg pivot_in_0_99;
     wire pivot_out_0_99;

     assign data_in_0_99 = data_in[DAT_W-100];

     always @(posedge clk) begin
        op_in_0_99 <= op_out_0_98;
        pivot_in_0_99 <= pivot_out_0_98;
        start_in_0_99 <= start_out_0_98;
        swap_in_0_99 <= swap_out_0_98;
     end
  
     processor_AB AB_0_99 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_99),
       .start_in   (start_in_0_99),
       .swap_in    (swap_in_0_99),
       .op_in      (op_in_0_99),
       .pivot_in   (pivot_in_0_99),
       .start_out  (start_out_0_99),
       .swap_out   (swap_out_0_99),
       .data_out   (data_out_0_99),
       .op_out     (op_out_0_99),
       .pivot_out  (pivot_out_0_99),
       .r          (r_0_99)
     );

  // row 0, col 100

     reg start_in_0_100;
     wire start_out_0_100;

     reg swap_in_0_100;
     wire swap_out_0_100;

     reg [1:0] op_in_0_100;
     wire [1:0] op_out_0_100;

     wire r_0_100;

     wire data_in_0_100;
     wire data_out_0_100;

     reg pivot_in_0_100;
     wire pivot_out_0_100;

     assign data_in_0_100 = data_in[DAT_W-101];

     always @(posedge clk) begin
        op_in_0_100 <= op_out_0_99;
        pivot_in_0_100 <= pivot_out_0_99;
        start_in_0_100 <= start_out_0_99;
        swap_in_0_100 <= swap_out_0_99;
     end
  
     processor_AB AB_0_100 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_100),
       .start_in   (start_in_0_100),
       .swap_in    (swap_in_0_100),
       .op_in      (op_in_0_100),
       .pivot_in   (pivot_in_0_100),
       .start_out  (start_out_0_100),
       .swap_out   (swap_out_0_100),
       .data_out   (data_out_0_100),
       .op_out     (op_out_0_100),
       .pivot_out  (pivot_out_0_100),
       .r          (r_0_100)
     );

  // row 0, col 101

     reg start_in_0_101;
     wire start_out_0_101;

     reg swap_in_0_101;
     wire swap_out_0_101;

     reg [1:0] op_in_0_101;
     wire [1:0] op_out_0_101;

     wire r_0_101;

     wire data_in_0_101;
     wire data_out_0_101;

     reg pivot_in_0_101;
     wire pivot_out_0_101;

     assign data_in_0_101 = data_in[DAT_W-102];

     always @(posedge clk) begin
        op_in_0_101 <= op_out_0_100;
        pivot_in_0_101 <= pivot_out_0_100;
        start_in_0_101 <= start_out_0_100;
        swap_in_0_101 <= swap_out_0_100;
     end
  
     processor_AB AB_0_101 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_101),
       .start_in   (start_in_0_101),
       .swap_in    (swap_in_0_101),
       .op_in      (op_in_0_101),
       .pivot_in   (pivot_in_0_101),
       .start_out  (start_out_0_101),
       .swap_out   (swap_out_0_101),
       .data_out   (data_out_0_101),
       .op_out     (op_out_0_101),
       .pivot_out  (pivot_out_0_101),
       .r          (r_0_101)
     );

  // row 0, col 102

     reg start_in_0_102;
     wire start_out_0_102;

     reg swap_in_0_102;
     wire swap_out_0_102;

     reg [1:0] op_in_0_102;
     wire [1:0] op_out_0_102;

     wire r_0_102;

     wire data_in_0_102;
     wire data_out_0_102;

     reg pivot_in_0_102;
     wire pivot_out_0_102;

     assign data_in_0_102 = data_in[DAT_W-103];

     always @(posedge clk) begin
        op_in_0_102 <= op_out_0_101;
        pivot_in_0_102 <= pivot_out_0_101;
        start_in_0_102 <= start_out_0_101;
        swap_in_0_102 <= swap_out_0_101;
     end
  
     processor_AB AB_0_102 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_102),
       .start_in   (start_in_0_102),
       .swap_in    (swap_in_0_102),
       .op_in      (op_in_0_102),
       .pivot_in   (pivot_in_0_102),
       .start_out  (start_out_0_102),
       .swap_out   (swap_out_0_102),
       .data_out   (data_out_0_102),
       .op_out     (op_out_0_102),
       .pivot_out  (pivot_out_0_102),
       .r          (r_0_102)
     );

  // row 0, col 103

     reg start_in_0_103;
     wire start_out_0_103;

     reg swap_in_0_103;
     wire swap_out_0_103;

     reg [1:0] op_in_0_103;
     wire [1:0] op_out_0_103;

     wire r_0_103;

     wire data_in_0_103;
     wire data_out_0_103;

     reg pivot_in_0_103;
     wire pivot_out_0_103;

     assign data_in_0_103 = data_in[DAT_W-104];

     always @(posedge clk) begin
        op_in_0_103 <= op_out_0_102;
        pivot_in_0_103 <= pivot_out_0_102;
        start_in_0_103 <= start_out_0_102;
        swap_in_0_103 <= swap_out_0_102;
     end
  
     processor_AB AB_0_103 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_103),
       .start_in   (start_in_0_103),
       .swap_in    (swap_in_0_103),
       .op_in      (op_in_0_103),
       .pivot_in   (pivot_in_0_103),
       .start_out  (start_out_0_103),
       .swap_out   (swap_out_0_103),
       .data_out   (data_out_0_103),
       .op_out     (op_out_0_103),
       .pivot_out  (pivot_out_0_103),
       .r          (r_0_103)
     );

  // row 0, col 104

     reg start_in_0_104;
     wire start_out_0_104;

     reg swap_in_0_104;
     wire swap_out_0_104;

     reg [1:0] op_in_0_104;
     wire [1:0] op_out_0_104;

     wire r_0_104;

     wire data_in_0_104;
     wire data_out_0_104;

     reg pivot_in_0_104;
     wire pivot_out_0_104;

     assign data_in_0_104 = data_in[DAT_W-105];

     always @(posedge clk) begin
        op_in_0_104 <= op_out_0_103;
        pivot_in_0_104 <= pivot_out_0_103;
        start_in_0_104 <= start_out_0_103;
        swap_in_0_104 <= swap_out_0_103;
     end
  
     processor_AB AB_0_104 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_104),
       .start_in   (start_in_0_104),
       .swap_in    (swap_in_0_104),
       .op_in      (op_in_0_104),
       .pivot_in   (pivot_in_0_104),
       .start_out  (start_out_0_104),
       .swap_out   (swap_out_0_104),
       .data_out   (data_out_0_104),
       .op_out     (op_out_0_104),
       .pivot_out  (pivot_out_0_104),
       .r          (r_0_104)
     );

  // row 0, col 105

     reg start_in_0_105;
     wire start_out_0_105;

     reg swap_in_0_105;
     wire swap_out_0_105;

     reg [1:0] op_in_0_105;
     wire [1:0] op_out_0_105;

     wire r_0_105;

     wire data_in_0_105;
     wire data_out_0_105;

     reg pivot_in_0_105;
     wire pivot_out_0_105;

     assign data_in_0_105 = data_in[DAT_W-106];

     always @(posedge clk) begin
        op_in_0_105 <= op_out_0_104;
        pivot_in_0_105 <= pivot_out_0_104;
        start_in_0_105 <= start_out_0_104;
        swap_in_0_105 <= swap_out_0_104;
     end
  
     processor_AB AB_0_105 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_105),
       .start_in   (start_in_0_105),
       .swap_in    (swap_in_0_105),
       .op_in      (op_in_0_105),
       .pivot_in   (pivot_in_0_105),
       .start_out  (start_out_0_105),
       .swap_out   (swap_out_0_105),
       .data_out   (data_out_0_105),
       .op_out     (op_out_0_105),
       .pivot_out  (pivot_out_0_105),
       .r          (r_0_105)
     );

  // row 0, col 106

     reg start_in_0_106;
     wire start_out_0_106;

     reg swap_in_0_106;
     wire swap_out_0_106;

     reg [1:0] op_in_0_106;
     wire [1:0] op_out_0_106;

     wire r_0_106;

     wire data_in_0_106;
     wire data_out_0_106;

     reg pivot_in_0_106;
     wire pivot_out_0_106;

     assign data_in_0_106 = data_in[DAT_W-107];

     always @(posedge clk) begin
        op_in_0_106 <= op_out_0_105;
        pivot_in_0_106 <= pivot_out_0_105;
        start_in_0_106 <= start_out_0_105;
        swap_in_0_106 <= swap_out_0_105;
     end
  
     processor_AB AB_0_106 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_106),
       .start_in   (start_in_0_106),
       .swap_in    (swap_in_0_106),
       .op_in      (op_in_0_106),
       .pivot_in   (pivot_in_0_106),
       .start_out  (start_out_0_106),
       .swap_out   (swap_out_0_106),
       .data_out   (data_out_0_106),
       .op_out     (op_out_0_106),
       .pivot_out  (pivot_out_0_106),
       .r          (r_0_106)
     );

  // row 0, col 107

     reg start_in_0_107;
     wire start_out_0_107;

     reg swap_in_0_107;
     wire swap_out_0_107;

     reg [1:0] op_in_0_107;
     wire [1:0] op_out_0_107;

     wire r_0_107;

     wire data_in_0_107;
     wire data_out_0_107;

     reg pivot_in_0_107;
     wire pivot_out_0_107;

     assign data_in_0_107 = data_in[DAT_W-108];

     always @(posedge clk) begin
        op_in_0_107 <= op_out_0_106;
        pivot_in_0_107 <= pivot_out_0_106;
        start_in_0_107 <= start_out_0_106;
        swap_in_0_107 <= swap_out_0_106;
     end
  
     processor_AB AB_0_107 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_107),
       .start_in   (start_in_0_107),
       .swap_in    (swap_in_0_107),
       .op_in      (op_in_0_107),
       .pivot_in   (pivot_in_0_107),
       .start_out  (start_out_0_107),
       .swap_out   (swap_out_0_107),
       .data_out   (data_out_0_107),
       .op_out     (op_out_0_107),
       .pivot_out  (pivot_out_0_107),
       .r          (r_0_107)
     );

  // row 0, col 108

     reg start_in_0_108;
     wire start_out_0_108;

     reg swap_in_0_108;
     wire swap_out_0_108;

     reg [1:0] op_in_0_108;
     wire [1:0] op_out_0_108;

     wire r_0_108;

     wire data_in_0_108;
     wire data_out_0_108;

     reg pivot_in_0_108;
     wire pivot_out_0_108;

     assign data_in_0_108 = data_in[DAT_W-109];

     always @(posedge clk) begin
        op_in_0_108 <= op_out_0_107;
        pivot_in_0_108 <= pivot_out_0_107;
        start_in_0_108 <= start_out_0_107;
        swap_in_0_108 <= swap_out_0_107;
     end
  
     processor_AB AB_0_108 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_108),
       .start_in   (start_in_0_108),
       .swap_in    (swap_in_0_108),
       .op_in      (op_in_0_108),
       .pivot_in   (pivot_in_0_108),
       .start_out  (start_out_0_108),
       .swap_out   (swap_out_0_108),
       .data_out   (data_out_0_108),
       .op_out     (op_out_0_108),
       .pivot_out  (pivot_out_0_108),
       .r          (r_0_108)
     );

  // row 0, col 109

     reg start_in_0_109;
     wire start_out_0_109;

     reg swap_in_0_109;
     wire swap_out_0_109;

     reg [1:0] op_in_0_109;
     wire [1:0] op_out_0_109;

     wire r_0_109;

     wire data_in_0_109;
     wire data_out_0_109;

     reg pivot_in_0_109;
     wire pivot_out_0_109;

     assign data_in_0_109 = data_in[DAT_W-110];

     always @(posedge clk) begin
        op_in_0_109 <= op_out_0_108;
        pivot_in_0_109 <= pivot_out_0_108;
        start_in_0_109 <= start_out_0_108;
        swap_in_0_109 <= swap_out_0_108;
     end
  
     processor_AB AB_0_109 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_109),
       .start_in   (start_in_0_109),
       .swap_in    (swap_in_0_109),
       .op_in      (op_in_0_109),
       .pivot_in   (pivot_in_0_109),
       .start_out  (start_out_0_109),
       .swap_out   (swap_out_0_109),
       .data_out   (data_out_0_109),
       .op_out     (op_out_0_109),
       .pivot_out  (pivot_out_0_109),
       .r          (r_0_109)
     );

  // row 0, col 110

     reg start_in_0_110;
     wire start_out_0_110;

     reg swap_in_0_110;
     wire swap_out_0_110;

     reg [1:0] op_in_0_110;
     wire [1:0] op_out_0_110;

     wire r_0_110;

     wire data_in_0_110;
     wire data_out_0_110;

     reg pivot_in_0_110;
     wire pivot_out_0_110;

     assign data_in_0_110 = data_in[DAT_W-111];

     always @(posedge clk) begin
        op_in_0_110 <= op_out_0_109;
        pivot_in_0_110 <= pivot_out_0_109;
        start_in_0_110 <= start_out_0_109;
        swap_in_0_110 <= swap_out_0_109;
     end
  
     processor_AB AB_0_110 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_110),
       .start_in   (start_in_0_110),
       .swap_in    (swap_in_0_110),
       .op_in      (op_in_0_110),
       .pivot_in   (pivot_in_0_110),
       .start_out  (start_out_0_110),
       .swap_out   (swap_out_0_110),
       .data_out   (data_out_0_110),
       .op_out     (op_out_0_110),
       .pivot_out  (pivot_out_0_110),
       .r          (r_0_110)
     );

  // row 0, col 111

     reg start_in_0_111;
     wire start_out_0_111;

     reg swap_in_0_111;
     wire swap_out_0_111;

     reg [1:0] op_in_0_111;
     wire [1:0] op_out_0_111;

     wire r_0_111;

     wire data_in_0_111;
     wire data_out_0_111;

     reg pivot_in_0_111;
     wire pivot_out_0_111;

     assign data_in_0_111 = data_in[DAT_W-112];

     always @(posedge clk) begin
        op_in_0_111 <= op_out_0_110;
        pivot_in_0_111 <= pivot_out_0_110;
        start_in_0_111 <= start_out_0_110;
        swap_in_0_111 <= swap_out_0_110;
     end
  
     processor_AB AB_0_111 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_111),
       .start_in   (start_in_0_111),
       .swap_in    (swap_in_0_111),
       .op_in      (op_in_0_111),
       .pivot_in   (pivot_in_0_111),
       .start_out  (start_out_0_111),
       .swap_out   (swap_out_0_111),
       .data_out   (data_out_0_111),
       .op_out     (op_out_0_111),
       .pivot_out  (pivot_out_0_111),
       .r          (r_0_111)
     );

  // row 0, col 112

     reg start_in_0_112;
     wire start_out_0_112;

     reg swap_in_0_112;
     wire swap_out_0_112;

     reg [1:0] op_in_0_112;
     wire [1:0] op_out_0_112;

     wire r_0_112;

     wire data_in_0_112;
     wire data_out_0_112;

     reg pivot_in_0_112;
     wire pivot_out_0_112;

     assign data_in_0_112 = data_in[DAT_W-113];

     always @(posedge clk) begin
        op_in_0_112 <= op_out_0_111;
        pivot_in_0_112 <= pivot_out_0_111;
        start_in_0_112 <= start_out_0_111;
        swap_in_0_112 <= swap_out_0_111;
     end
  
     processor_AB AB_0_112 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_112),
       .start_in   (start_in_0_112),
       .swap_in    (swap_in_0_112),
       .op_in      (op_in_0_112),
       .pivot_in   (pivot_in_0_112),
       .start_out  (start_out_0_112),
       .swap_out   (swap_out_0_112),
       .data_out   (data_out_0_112),
       .op_out     (op_out_0_112),
       .pivot_out  (pivot_out_0_112),
       .r          (r_0_112)
     );

  // row 0, col 113

     reg start_in_0_113;
     wire start_out_0_113;

     reg swap_in_0_113;
     wire swap_out_0_113;

     reg [1:0] op_in_0_113;
     wire [1:0] op_out_0_113;

     wire r_0_113;

     wire data_in_0_113;
     wire data_out_0_113;

     reg pivot_in_0_113;
     wire pivot_out_0_113;

     assign data_in_0_113 = data_in[DAT_W-114];

     always @(posedge clk) begin
        op_in_0_113 <= op_out_0_112;
        pivot_in_0_113 <= pivot_out_0_112;
        start_in_0_113 <= start_out_0_112;
        swap_in_0_113 <= swap_out_0_112;
     end
  
     processor_AB AB_0_113 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_113),
       .start_in   (start_in_0_113),
       .swap_in    (swap_in_0_113),
       .op_in      (op_in_0_113),
       .pivot_in   (pivot_in_0_113),
       .start_out  (start_out_0_113),
       .swap_out   (swap_out_0_113),
       .data_out   (data_out_0_113),
       .op_out     (op_out_0_113),
       .pivot_out  (pivot_out_0_113),
       .r          (r_0_113)
     );

  // row 0, col 114

     reg start_in_0_114;
     wire start_out_0_114;

     reg swap_in_0_114;
     wire swap_out_0_114;

     reg [1:0] op_in_0_114;
     wire [1:0] op_out_0_114;

     wire r_0_114;

     wire data_in_0_114;
     wire data_out_0_114;

     reg pivot_in_0_114;
     wire pivot_out_0_114;

     assign data_in_0_114 = data_in[DAT_W-115];

     always @(posedge clk) begin
        op_in_0_114 <= op_out_0_113;
        pivot_in_0_114 <= pivot_out_0_113;
        start_in_0_114 <= start_out_0_113;
        swap_in_0_114 <= swap_out_0_113;
     end
  
     processor_AB AB_0_114 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_114),
       .start_in   (start_in_0_114),
       .swap_in    (swap_in_0_114),
       .op_in      (op_in_0_114),
       .pivot_in   (pivot_in_0_114),
       .start_out  (start_out_0_114),
       .swap_out   (swap_out_0_114),
       .data_out   (data_out_0_114),
       .op_out     (op_out_0_114),
       .pivot_out  (pivot_out_0_114),
       .r          (r_0_114)
     );

  // row 0, col 115

     reg start_in_0_115;
     wire start_out_0_115;

     reg swap_in_0_115;
     wire swap_out_0_115;

     reg [1:0] op_in_0_115;
     wire [1:0] op_out_0_115;

     wire r_0_115;

     wire data_in_0_115;
     wire data_out_0_115;

     reg pivot_in_0_115;
     wire pivot_out_0_115;

     assign data_in_0_115 = data_in[DAT_W-116];

     always @(posedge clk) begin
        op_in_0_115 <= op_out_0_114;
        pivot_in_0_115 <= pivot_out_0_114;
        start_in_0_115 <= start_out_0_114;
        swap_in_0_115 <= swap_out_0_114;
     end
  
     processor_AB AB_0_115 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_115),
       .start_in   (start_in_0_115),
       .swap_in    (swap_in_0_115),
       .op_in      (op_in_0_115),
       .pivot_in   (pivot_in_0_115),
       .start_out  (start_out_0_115),
       .swap_out   (swap_out_0_115),
       .data_out   (data_out_0_115),
       .op_out     (op_out_0_115),
       .pivot_out  (pivot_out_0_115),
       .r          (r_0_115)
     );

  // row 0, col 116

     reg start_in_0_116;
     wire start_out_0_116;

     reg swap_in_0_116;
     wire swap_out_0_116;

     reg [1:0] op_in_0_116;
     wire [1:0] op_out_0_116;

     wire r_0_116;

     wire data_in_0_116;
     wire data_out_0_116;

     reg pivot_in_0_116;
     wire pivot_out_0_116;

     assign data_in_0_116 = data_in[DAT_W-117];

     always @(posedge clk) begin
        op_in_0_116 <= op_out_0_115;
        pivot_in_0_116 <= pivot_out_0_115;
        start_in_0_116 <= start_out_0_115;
        swap_in_0_116 <= swap_out_0_115;
     end
  
     processor_AB AB_0_116 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_116),
       .start_in   (start_in_0_116),
       .swap_in    (swap_in_0_116),
       .op_in      (op_in_0_116),
       .pivot_in   (pivot_in_0_116),
       .start_out  (start_out_0_116),
       .swap_out   (swap_out_0_116),
       .data_out   (data_out_0_116),
       .op_out     (op_out_0_116),
       .pivot_out  (pivot_out_0_116),
       .r          (r_0_116)
     );

  // row 0, col 117

     reg start_in_0_117;
     wire start_out_0_117;

     reg swap_in_0_117;
     wire swap_out_0_117;

     reg [1:0] op_in_0_117;
     wire [1:0] op_out_0_117;

     wire r_0_117;

     wire data_in_0_117;
     wire data_out_0_117;

     reg pivot_in_0_117;
     wire pivot_out_0_117;

     assign data_in_0_117 = data_in[DAT_W-118];

     always @(posedge clk) begin
        op_in_0_117 <= op_out_0_116;
        pivot_in_0_117 <= pivot_out_0_116;
        start_in_0_117 <= start_out_0_116;
        swap_in_0_117 <= swap_out_0_116;
     end
  
     processor_AB AB_0_117 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_117),
       .start_in   (start_in_0_117),
       .swap_in    (swap_in_0_117),
       .op_in      (op_in_0_117),
       .pivot_in   (pivot_in_0_117),
       .start_out  (start_out_0_117),
       .swap_out   (swap_out_0_117),
       .data_out   (data_out_0_117),
       .op_out     (op_out_0_117),
       .pivot_out  (pivot_out_0_117),
       .r          (r_0_117)
     );

  // row 0, col 118

     reg start_in_0_118;
     wire start_out_0_118;

     reg swap_in_0_118;
     wire swap_out_0_118;

     reg [1:0] op_in_0_118;
     wire [1:0] op_out_0_118;

     wire r_0_118;

     wire data_in_0_118;
     wire data_out_0_118;

     reg pivot_in_0_118;
     wire pivot_out_0_118;

     assign data_in_0_118 = data_in[DAT_W-119];

     always @(posedge clk) begin
        op_in_0_118 <= op_out_0_117;
        pivot_in_0_118 <= pivot_out_0_117;
        start_in_0_118 <= start_out_0_117;
        swap_in_0_118 <= swap_out_0_117;
     end
  
     processor_AB AB_0_118 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_118),
       .start_in   (start_in_0_118),
       .swap_in    (swap_in_0_118),
       .op_in      (op_in_0_118),
       .pivot_in   (pivot_in_0_118),
       .start_out  (start_out_0_118),
       .swap_out   (swap_out_0_118),
       .data_out   (data_out_0_118),
       .op_out     (op_out_0_118),
       .pivot_out  (pivot_out_0_118),
       .r          (r_0_118)
     );

  // row 0, col 119

     reg start_in_0_119;
     wire start_out_0_119;

     reg swap_in_0_119;
     wire swap_out_0_119;

     reg [1:0] op_in_0_119;
     wire [1:0] op_out_0_119;

     wire r_0_119;

     wire data_in_0_119;
     wire data_out_0_119;

     reg pivot_in_0_119;
     wire pivot_out_0_119;

     assign data_in_0_119 = data_in[DAT_W-120];

     always @(posedge clk) begin
        op_in_0_119 <= op_out_0_118;
        pivot_in_0_119 <= pivot_out_0_118;
        start_in_0_119 <= start_out_0_118;
        swap_in_0_119 <= swap_out_0_118;
     end
  
     processor_AB AB_0_119 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_119),
       .start_in   (start_in_0_119),
       .swap_in    (swap_in_0_119),
       .op_in      (op_in_0_119),
       .pivot_in   (pivot_in_0_119),
       .start_out  (start_out_0_119),
       .swap_out   (swap_out_0_119),
       .data_out   (data_out_0_119),
       .op_out     (op_out_0_119),
       .pivot_out  (pivot_out_0_119),
       .r          (r_0_119)
     );

  // row 0, col 120

     reg start_in_0_120;
     wire start_out_0_120;

     reg swap_in_0_120;
     wire swap_out_0_120;

     reg [1:0] op_in_0_120;
     wire [1:0] op_out_0_120;

     wire r_0_120;

     wire data_in_0_120;
     wire data_out_0_120;

     reg pivot_in_0_120;
     wire pivot_out_0_120;

     assign data_in_0_120 = data_in[DAT_W-121];

     always @(posedge clk) begin
        op_in_0_120 <= op_out_0_119;
        pivot_in_0_120 <= pivot_out_0_119;
        start_in_0_120 <= start_out_0_119;
        swap_in_0_120 <= swap_out_0_119;
     end
  
     processor_AB AB_0_120 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_120),
       .start_in   (start_in_0_120),
       .swap_in    (swap_in_0_120),
       .op_in      (op_in_0_120),
       .pivot_in   (pivot_in_0_120),
       .start_out  (start_out_0_120),
       .swap_out   (swap_out_0_120),
       .data_out   (data_out_0_120),
       .op_out     (op_out_0_120),
       .pivot_out  (pivot_out_0_120),
       .r          (r_0_120)
     );

  // row 0, col 121

     reg start_in_0_121;
     wire start_out_0_121;

     reg swap_in_0_121;
     wire swap_out_0_121;

     reg [1:0] op_in_0_121;
     wire [1:0] op_out_0_121;

     wire r_0_121;

     wire data_in_0_121;
     wire data_out_0_121;

     reg pivot_in_0_121;
     wire pivot_out_0_121;

     assign data_in_0_121 = data_in[DAT_W-122];

     always @(posedge clk) begin
        op_in_0_121 <= op_out_0_120;
        pivot_in_0_121 <= pivot_out_0_120;
        start_in_0_121 <= start_out_0_120;
        swap_in_0_121 <= swap_out_0_120;
     end
  
     processor_AB AB_0_121 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_121),
       .start_in   (start_in_0_121),
       .swap_in    (swap_in_0_121),
       .op_in      (op_in_0_121),
       .pivot_in   (pivot_in_0_121),
       .start_out  (start_out_0_121),
       .swap_out   (swap_out_0_121),
       .data_out   (data_out_0_121),
       .op_out     (op_out_0_121),
       .pivot_out  (pivot_out_0_121),
       .r          (r_0_121)
     );

  // row 0, col 122

     reg start_in_0_122;
     wire start_out_0_122;

     reg swap_in_0_122;
     wire swap_out_0_122;

     reg [1:0] op_in_0_122;
     wire [1:0] op_out_0_122;

     wire r_0_122;

     wire data_in_0_122;
     wire data_out_0_122;

     reg pivot_in_0_122;
     wire pivot_out_0_122;

     assign data_in_0_122 = data_in[DAT_W-123];

     always @(posedge clk) begin
        op_in_0_122 <= op_out_0_121;
        pivot_in_0_122 <= pivot_out_0_121;
        start_in_0_122 <= start_out_0_121;
        swap_in_0_122 <= swap_out_0_121;
     end
  
     processor_AB AB_0_122 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_122),
       .start_in   (start_in_0_122),
       .swap_in    (swap_in_0_122),
       .op_in      (op_in_0_122),
       .pivot_in   (pivot_in_0_122),
       .start_out  (start_out_0_122),
       .swap_out   (swap_out_0_122),
       .data_out   (data_out_0_122),
       .op_out     (op_out_0_122),
       .pivot_out  (pivot_out_0_122),
       .r          (r_0_122)
     );

  // row 0, col 123

     reg start_in_0_123;
     wire start_out_0_123;

     reg swap_in_0_123;
     wire swap_out_0_123;

     reg [1:0] op_in_0_123;
     wire [1:0] op_out_0_123;

     wire r_0_123;

     wire data_in_0_123;
     wire data_out_0_123;

     reg pivot_in_0_123;
     wire pivot_out_0_123;

     assign data_in_0_123 = data_in[DAT_W-124];

     always @(posedge clk) begin
        op_in_0_123 <= op_out_0_122;
        pivot_in_0_123 <= pivot_out_0_122;
        start_in_0_123 <= start_out_0_122;
        swap_in_0_123 <= swap_out_0_122;
     end
  
     processor_AB AB_0_123 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_123),
       .start_in   (start_in_0_123),
       .swap_in    (swap_in_0_123),
       .op_in      (op_in_0_123),
       .pivot_in   (pivot_in_0_123),
       .start_out  (start_out_0_123),
       .swap_out   (swap_out_0_123),
       .data_out   (data_out_0_123),
       .op_out     (op_out_0_123),
       .pivot_out  (pivot_out_0_123),
       .r          (r_0_123)
     );

  // row 0, col 124

     reg start_in_0_124;
     wire start_out_0_124;

     reg swap_in_0_124;
     wire swap_out_0_124;

     reg [1:0] op_in_0_124;
     wire [1:0] op_out_0_124;

     wire r_0_124;

     wire data_in_0_124;
     wire data_out_0_124;

     reg pivot_in_0_124;
     wire pivot_out_0_124;

     assign data_in_0_124 = data_in[DAT_W-125];

     always @(posedge clk) begin
        op_in_0_124 <= op_out_0_123;
        pivot_in_0_124 <= pivot_out_0_123;
        start_in_0_124 <= start_out_0_123;
        swap_in_0_124 <= swap_out_0_123;
     end
  
     processor_AB AB_0_124 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_124),
       .start_in   (start_in_0_124),
       .swap_in    (swap_in_0_124),
       .op_in      (op_in_0_124),
       .pivot_in   (pivot_in_0_124),
       .start_out  (start_out_0_124),
       .swap_out   (swap_out_0_124),
       .data_out   (data_out_0_124),
       .op_out     (op_out_0_124),
       .pivot_out  (pivot_out_0_124),
       .r          (r_0_124)
     );

  // row 0, col 125

     reg start_in_0_125;
     wire start_out_0_125;

     reg swap_in_0_125;
     wire swap_out_0_125;

     reg [1:0] op_in_0_125;
     wire [1:0] op_out_0_125;

     wire r_0_125;

     wire data_in_0_125;
     wire data_out_0_125;

     reg pivot_in_0_125;
     wire pivot_out_0_125;

     assign data_in_0_125 = data_in[DAT_W-126];

     always @(posedge clk) begin
        op_in_0_125 <= op_out_0_124;
        pivot_in_0_125 <= pivot_out_0_124;
        start_in_0_125 <= start_out_0_124;
        swap_in_0_125 <= swap_out_0_124;
     end
  
     processor_AB AB_0_125 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_125),
       .start_in   (start_in_0_125),
       .swap_in    (swap_in_0_125),
       .op_in      (op_in_0_125),
       .pivot_in   (pivot_in_0_125),
       .start_out  (start_out_0_125),
       .swap_out   (swap_out_0_125),
       .data_out   (data_out_0_125),
       .op_out     (op_out_0_125),
       .pivot_out  (pivot_out_0_125),
       .r          (r_0_125)
     );

  // row 0, col 126

     reg start_in_0_126;
     wire start_out_0_126;

     reg swap_in_0_126;
     wire swap_out_0_126;

     reg [1:0] op_in_0_126;
     wire [1:0] op_out_0_126;

     wire r_0_126;

     wire data_in_0_126;
     wire data_out_0_126;

     reg pivot_in_0_126;
     wire pivot_out_0_126;

     assign data_in_0_126 = data_in[DAT_W-127];

     always @(posedge clk) begin
        op_in_0_126 <= op_out_0_125;
        pivot_in_0_126 <= pivot_out_0_125;
        start_in_0_126 <= start_out_0_125;
        swap_in_0_126 <= swap_out_0_125;
     end
  
     processor_AB AB_0_126 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_126),
       .start_in   (start_in_0_126),
       .swap_in    (swap_in_0_126),
       .op_in      (op_in_0_126),
       .pivot_in   (pivot_in_0_126),
       .start_out  (start_out_0_126),
       .swap_out   (swap_out_0_126),
       .data_out   (data_out_0_126),
       .op_out     (op_out_0_126),
       .pivot_out  (pivot_out_0_126),
       .r          (r_0_126)
     );

  // row 0, col 127

     reg start_in_0_127;
     wire start_out_0_127;

     reg swap_in_0_127;
     wire swap_out_0_127;

     reg [1:0] op_in_0_127;
     wire [1:0] op_out_0_127;

     wire r_0_127;

     wire data_in_0_127;
     wire data_out_0_127;

     reg pivot_in_0_127;
     wire pivot_out_0_127;

     assign data_in_0_127 = data_in[DAT_W-128];

     always @(posedge clk) begin
        op_in_0_127 <= op_out_0_126;
        pivot_in_0_127 <= pivot_out_0_126;
        start_in_0_127 <= start_out_0_126;
        swap_in_0_127 <= swap_out_0_126;
     end
  
     processor_AB AB_0_127 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_127),
       .start_in   (start_in_0_127),
       .swap_in    (swap_in_0_127),
       .op_in      (op_in_0_127),
       .pivot_in   (pivot_in_0_127),
       .start_out  (start_out_0_127),
       .swap_out   (swap_out_0_127),
       .data_out   (data_out_0_127),
       .op_out     (op_out_0_127),
       .pivot_out  (pivot_out_0_127),
       .r          (r_0_127)
     );

  // row 0, col 128

     reg start_in_0_128;
     wire start_out_0_128;

     reg swap_in_0_128;
     wire swap_out_0_128;

     reg [1:0] op_in_0_128;
     wire [1:0] op_out_0_128;

     wire r_0_128;

     wire data_in_0_128;
     wire data_out_0_128;

     reg pivot_in_0_128;
     wire pivot_out_0_128;

     assign data_in_0_128 = data_in[DAT_W-129];

     always @(posedge clk) begin
        op_in_0_128 <= op_out_0_127;
        pivot_in_0_128 <= pivot_out_0_127;
        start_in_0_128 <= start_out_0_127;
        swap_in_0_128 <= swap_out_0_127;
     end
  
     processor_AB AB_0_128 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_128),
       .start_in   (start_in_0_128),
       .swap_in    (swap_in_0_128),
       .op_in      (op_in_0_128),
       .pivot_in   (pivot_in_0_128),
       .start_out  (start_out_0_128),
       .swap_out   (swap_out_0_128),
       .data_out   (data_out_0_128),
       .op_out     (op_out_0_128),
       .pivot_out  (pivot_out_0_128),
       .r          (r_0_128)
     );

  // row 0, col 129

     reg start_in_0_129;
     wire start_out_0_129;

     reg swap_in_0_129;
     wire swap_out_0_129;

     reg [1:0] op_in_0_129;
     wire [1:0] op_out_0_129;

     wire r_0_129;

     wire data_in_0_129;
     wire data_out_0_129;

     reg pivot_in_0_129;
     wire pivot_out_0_129;

     assign data_in_0_129 = data_in[DAT_W-130];

     always @(posedge clk) begin
        op_in_0_129 <= op_out_0_128;
        pivot_in_0_129 <= pivot_out_0_128;
        start_in_0_129 <= start_out_0_128;
        swap_in_0_129 <= swap_out_0_128;
     end
  
     processor_AB AB_0_129 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_129),
       .start_in   (start_in_0_129),
       .swap_in    (swap_in_0_129),
       .op_in      (op_in_0_129),
       .pivot_in   (pivot_in_0_129),
       .start_out  (start_out_0_129),
       .swap_out   (swap_out_0_129),
       .data_out   (data_out_0_129),
       .op_out     (op_out_0_129),
       .pivot_out  (pivot_out_0_129),
       .r          (r_0_129)
     );

  // row 0, col 130

     reg start_in_0_130;
     wire start_out_0_130;

     reg swap_in_0_130;
     wire swap_out_0_130;

     reg [1:0] op_in_0_130;
     wire [1:0] op_out_0_130;

     wire r_0_130;

     wire data_in_0_130;
     wire data_out_0_130;

     reg pivot_in_0_130;
     wire pivot_out_0_130;

     assign data_in_0_130 = data_in[DAT_W-131];

     always @(posedge clk) begin
        op_in_0_130 <= op_out_0_129;
        pivot_in_0_130 <= pivot_out_0_129;
        start_in_0_130 <= start_out_0_129;
        swap_in_0_130 <= swap_out_0_129;
     end
  
     processor_AB AB_0_130 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_130),
       .start_in   (start_in_0_130),
       .swap_in    (swap_in_0_130),
       .op_in      (op_in_0_130),
       .pivot_in   (pivot_in_0_130),
       .start_out  (start_out_0_130),
       .swap_out   (swap_out_0_130),
       .data_out   (data_out_0_130),
       .op_out     (op_out_0_130),
       .pivot_out  (pivot_out_0_130),
       .r          (r_0_130)
     );

  // row 0, col 131

     reg start_in_0_131;
     wire start_out_0_131;

     reg swap_in_0_131;
     wire swap_out_0_131;

     reg [1:0] op_in_0_131;
     wire [1:0] op_out_0_131;

     wire r_0_131;

     wire data_in_0_131;
     wire data_out_0_131;

     reg pivot_in_0_131;
     wire pivot_out_0_131;

     assign data_in_0_131 = data_in[DAT_W-132];

     always @(posedge clk) begin
        op_in_0_131 <= op_out_0_130;
        pivot_in_0_131 <= pivot_out_0_130;
        start_in_0_131 <= start_out_0_130;
        swap_in_0_131 <= swap_out_0_130;
     end
  
     processor_AB AB_0_131 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_131),
       .start_in   (start_in_0_131),
       .swap_in    (swap_in_0_131),
       .op_in      (op_in_0_131),
       .pivot_in   (pivot_in_0_131),
       .start_out  (start_out_0_131),
       .swap_out   (swap_out_0_131),
       .data_out   (data_out_0_131),
       .op_out     (op_out_0_131),
       .pivot_out  (pivot_out_0_131),
       .r          (r_0_131)
     );

  // row 0, col 132

     reg start_in_0_132;
     wire start_out_0_132;

     reg swap_in_0_132;
     wire swap_out_0_132;

     reg [1:0] op_in_0_132;
     wire [1:0] op_out_0_132;

     wire r_0_132;

     wire data_in_0_132;
     wire data_out_0_132;

     reg pivot_in_0_132;
     wire pivot_out_0_132;

     assign data_in_0_132 = data_in[DAT_W-133];

     always @(posedge clk) begin
        op_in_0_132 <= op_out_0_131;
        pivot_in_0_132 <= pivot_out_0_131;
        start_in_0_132 <= start_out_0_131;
        swap_in_0_132 <= swap_out_0_131;
     end
  
     processor_AB AB_0_132 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_132),
       .start_in   (start_in_0_132),
       .swap_in    (swap_in_0_132),
       .op_in      (op_in_0_132),
       .pivot_in   (pivot_in_0_132),
       .start_out  (start_out_0_132),
       .swap_out   (swap_out_0_132),
       .data_out   (data_out_0_132),
       .op_out     (op_out_0_132),
       .pivot_out  (pivot_out_0_132),
       .r          (r_0_132)
     );

  // row 0, col 133

     reg start_in_0_133;
     wire start_out_0_133;

     reg swap_in_0_133;
     wire swap_out_0_133;

     reg [1:0] op_in_0_133;
     wire [1:0] op_out_0_133;

     wire r_0_133;

     wire data_in_0_133;
     wire data_out_0_133;

     reg pivot_in_0_133;
     wire pivot_out_0_133;

     assign data_in_0_133 = data_in[DAT_W-134];

     always @(posedge clk) begin
        op_in_0_133 <= op_out_0_132;
        pivot_in_0_133 <= pivot_out_0_132;
        start_in_0_133 <= start_out_0_132;
        swap_in_0_133 <= swap_out_0_132;
     end
  
     processor_AB AB_0_133 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_133),
       .start_in   (start_in_0_133),
       .swap_in    (swap_in_0_133),
       .op_in      (op_in_0_133),
       .pivot_in   (pivot_in_0_133),
       .start_out  (start_out_0_133),
       .swap_out   (swap_out_0_133),
       .data_out   (data_out_0_133),
       .op_out     (op_out_0_133),
       .pivot_out  (pivot_out_0_133),
       .r          (r_0_133)
     );

  // row 0, col 134

     reg start_in_0_134;
     wire start_out_0_134;

     reg swap_in_0_134;
     wire swap_out_0_134;

     reg [1:0] op_in_0_134;
     wire [1:0] op_out_0_134;

     wire r_0_134;

     wire data_in_0_134;
     wire data_out_0_134;

     reg pivot_in_0_134;
     wire pivot_out_0_134;

     assign data_in_0_134 = data_in[DAT_W-135];

     always @(posedge clk) begin
        op_in_0_134 <= op_out_0_133;
        pivot_in_0_134 <= pivot_out_0_133;
        start_in_0_134 <= start_out_0_133;
        swap_in_0_134 <= swap_out_0_133;
     end
  
     processor_AB AB_0_134 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_134),
       .start_in   (start_in_0_134),
       .swap_in    (swap_in_0_134),
       .op_in      (op_in_0_134),
       .pivot_in   (pivot_in_0_134),
       .start_out  (start_out_0_134),
       .swap_out   (swap_out_0_134),
       .data_out   (data_out_0_134),
       .op_out     (op_out_0_134),
       .pivot_out  (pivot_out_0_134),
       .r          (r_0_134)
     );

  // row 0, col 135

     reg start_in_0_135;
     wire start_out_0_135;

     reg swap_in_0_135;
     wire swap_out_0_135;

     reg [1:0] op_in_0_135;
     wire [1:0] op_out_0_135;

     wire r_0_135;

     wire data_in_0_135;
     wire data_out_0_135;

     reg pivot_in_0_135;
     wire pivot_out_0_135;

     assign data_in_0_135 = data_in[DAT_W-136];

     always @(posedge clk) begin
        op_in_0_135 <= op_out_0_134;
        pivot_in_0_135 <= pivot_out_0_134;
        start_in_0_135 <= start_out_0_134;
        swap_in_0_135 <= swap_out_0_134;
     end
  
     processor_AB AB_0_135 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_135),
       .start_in   (start_in_0_135),
       .swap_in    (swap_in_0_135),
       .op_in      (op_in_0_135),
       .pivot_in   (pivot_in_0_135),
       .start_out  (start_out_0_135),
       .swap_out   (swap_out_0_135),
       .data_out   (data_out_0_135),
       .op_out     (op_out_0_135),
       .pivot_out  (pivot_out_0_135),
       .r          (r_0_135)
     );

  // row 0, col 136

     reg start_in_0_136;
     wire start_out_0_136;

     reg swap_in_0_136;
     wire swap_out_0_136;

     reg [1:0] op_in_0_136;
     wire [1:0] op_out_0_136;

     wire r_0_136;

     wire data_in_0_136;
     wire data_out_0_136;

     reg pivot_in_0_136;
     wire pivot_out_0_136;

     assign data_in_0_136 = data_in[DAT_W-137];

     always @(posedge clk) begin
        op_in_0_136 <= op_out_0_135;
        pivot_in_0_136 <= pivot_out_0_135;
        start_in_0_136 <= start_out_0_135;
        swap_in_0_136 <= swap_out_0_135;
     end
  
     processor_AB AB_0_136 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_136),
       .start_in   (start_in_0_136),
       .swap_in    (swap_in_0_136),
       .op_in      (op_in_0_136),
       .pivot_in   (pivot_in_0_136),
       .start_out  (start_out_0_136),
       .swap_out   (swap_out_0_136),
       .data_out   (data_out_0_136),
       .op_out     (op_out_0_136),
       .pivot_out  (pivot_out_0_136),
       .r          (r_0_136)
     );

  // row 0, col 137

     reg start_in_0_137;
     wire start_out_0_137;

     reg swap_in_0_137;
     wire swap_out_0_137;

     reg [1:0] op_in_0_137;
     wire [1:0] op_out_0_137;

     wire r_0_137;

     wire data_in_0_137;
     wire data_out_0_137;

     reg pivot_in_0_137;
     wire pivot_out_0_137;

     assign data_in_0_137 = data_in[DAT_W-138];

     always @(posedge clk) begin
        op_in_0_137 <= op_out_0_136;
        pivot_in_0_137 <= pivot_out_0_136;
        start_in_0_137 <= start_out_0_136;
        swap_in_0_137 <= swap_out_0_136;
     end
  
     processor_AB AB_0_137 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_137),
       .start_in   (start_in_0_137),
       .swap_in    (swap_in_0_137),
       .op_in      (op_in_0_137),
       .pivot_in   (pivot_in_0_137),
       .start_out  (start_out_0_137),
       .swap_out   (swap_out_0_137),
       .data_out   (data_out_0_137),
       .op_out     (op_out_0_137),
       .pivot_out  (pivot_out_0_137),
       .r          (r_0_137)
     );

  // row 0, col 138

     reg start_in_0_138;
     wire start_out_0_138;

     reg swap_in_0_138;
     wire swap_out_0_138;

     reg [1:0] op_in_0_138;
     wire [1:0] op_out_0_138;

     wire r_0_138;

     wire data_in_0_138;
     wire data_out_0_138;

     reg pivot_in_0_138;
     wire pivot_out_0_138;

     assign data_in_0_138 = data_in[DAT_W-139];

     always @(posedge clk) begin
        op_in_0_138 <= op_out_0_137;
        pivot_in_0_138 <= pivot_out_0_137;
        start_in_0_138 <= start_out_0_137;
        swap_in_0_138 <= swap_out_0_137;
     end
  
     processor_AB AB_0_138 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_138),
       .start_in   (start_in_0_138),
       .swap_in    (swap_in_0_138),
       .op_in      (op_in_0_138),
       .pivot_in   (pivot_in_0_138),
       .start_out  (start_out_0_138),
       .swap_out   (swap_out_0_138),
       .data_out   (data_out_0_138),
       .op_out     (op_out_0_138),
       .pivot_out  (pivot_out_0_138),
       .r          (r_0_138)
     );

  // row 0, col 139

     reg start_in_0_139;
     wire start_out_0_139;

     reg swap_in_0_139;
     wire swap_out_0_139;

     reg [1:0] op_in_0_139;
     wire [1:0] op_out_0_139;

     wire r_0_139;

     wire data_in_0_139;
     wire data_out_0_139;

     reg pivot_in_0_139;
     wire pivot_out_0_139;

     assign data_in_0_139 = data_in[DAT_W-140];

     always @(posedge clk) begin
        op_in_0_139 <= op_out_0_138;
        pivot_in_0_139 <= pivot_out_0_138;
        start_in_0_139 <= start_out_0_138;
        swap_in_0_139 <= swap_out_0_138;
     end
  
     processor_AB AB_0_139 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_139),
       .start_in   (start_in_0_139),
       .swap_in    (swap_in_0_139),
       .op_in      (op_in_0_139),
       .pivot_in   (pivot_in_0_139),
       .start_out  (start_out_0_139),
       .swap_out   (swap_out_0_139),
       .data_out   (data_out_0_139),
       .op_out     (op_out_0_139),
       .pivot_out  (pivot_out_0_139),
       .r          (r_0_139)
     );

  // row 0, col 140

     reg start_in_0_140;
     wire start_out_0_140;

     reg swap_in_0_140;
     wire swap_out_0_140;

     reg [1:0] op_in_0_140;
     wire [1:0] op_out_0_140;

     wire r_0_140;

     wire data_in_0_140;
     wire data_out_0_140;

     reg pivot_in_0_140;
     wire pivot_out_0_140;

     assign data_in_0_140 = data_in[DAT_W-141];

     always @(posedge clk) begin
        op_in_0_140 <= op_out_0_139;
        pivot_in_0_140 <= pivot_out_0_139;
        start_in_0_140 <= start_out_0_139;
        swap_in_0_140 <= swap_out_0_139;
     end
  
     processor_AB AB_0_140 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_140),
       .start_in   (start_in_0_140),
       .swap_in    (swap_in_0_140),
       .op_in      (op_in_0_140),
       .pivot_in   (pivot_in_0_140),
       .start_out  (start_out_0_140),
       .swap_out   (swap_out_0_140),
       .data_out   (data_out_0_140),
       .op_out     (op_out_0_140),
       .pivot_out  (pivot_out_0_140),
       .r          (r_0_140)
     );

  // row 0, col 141

     reg start_in_0_141;
     wire start_out_0_141;

     reg swap_in_0_141;
     wire swap_out_0_141;

     reg [1:0] op_in_0_141;
     wire [1:0] op_out_0_141;

     wire r_0_141;

     wire data_in_0_141;
     wire data_out_0_141;

     reg pivot_in_0_141;
     wire pivot_out_0_141;

     assign data_in_0_141 = data_in[DAT_W-142];

     always @(posedge clk) begin
        op_in_0_141 <= op_out_0_140;
        pivot_in_0_141 <= pivot_out_0_140;
        start_in_0_141 <= start_out_0_140;
        swap_in_0_141 <= swap_out_0_140;
     end
  
     processor_AB AB_0_141 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_141),
       .start_in   (start_in_0_141),
       .swap_in    (swap_in_0_141),
       .op_in      (op_in_0_141),
       .pivot_in   (pivot_in_0_141),
       .start_out  (start_out_0_141),
       .swap_out   (swap_out_0_141),
       .data_out   (data_out_0_141),
       .op_out     (op_out_0_141),
       .pivot_out  (pivot_out_0_141),
       .r          (r_0_141)
     );

  // row 0, col 142

     reg start_in_0_142;
     wire start_out_0_142;

     reg swap_in_0_142;
     wire swap_out_0_142;

     reg [1:0] op_in_0_142;
     wire [1:0] op_out_0_142;

     wire r_0_142;

     wire data_in_0_142;
     wire data_out_0_142;

     reg pivot_in_0_142;
     wire pivot_out_0_142;

     assign data_in_0_142 = data_in[DAT_W-143];

     always @(posedge clk) begin
        op_in_0_142 <= op_out_0_141;
        pivot_in_0_142 <= pivot_out_0_141;
        start_in_0_142 <= start_out_0_141;
        swap_in_0_142 <= swap_out_0_141;
     end
  
     processor_AB AB_0_142 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_142),
       .start_in   (start_in_0_142),
       .swap_in    (swap_in_0_142),
       .op_in      (op_in_0_142),
       .pivot_in   (pivot_in_0_142),
       .start_out  (start_out_0_142),
       .swap_out   (swap_out_0_142),
       .data_out   (data_out_0_142),
       .op_out     (op_out_0_142),
       .pivot_out  (pivot_out_0_142),
       .r          (r_0_142)
     );

  // row 0, col 143

     reg start_in_0_143;
     wire start_out_0_143;

     reg swap_in_0_143;
     wire swap_out_0_143;

     reg [1:0] op_in_0_143;
     wire [1:0] op_out_0_143;

     wire r_0_143;

     wire data_in_0_143;
     wire data_out_0_143;

     reg pivot_in_0_143;
     wire pivot_out_0_143;

     assign data_in_0_143 = data_in[DAT_W-144];

     always @(posedge clk) begin
        op_in_0_143 <= op_out_0_142;
        pivot_in_0_143 <= pivot_out_0_142;
        start_in_0_143 <= start_out_0_142;
        swap_in_0_143 <= swap_out_0_142;
     end
  
     processor_AB AB_0_143 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_143),
       .start_in   (start_in_0_143),
       .swap_in    (swap_in_0_143),
       .op_in      (op_in_0_143),
       .pivot_in   (pivot_in_0_143),
       .start_out  (start_out_0_143),
       .swap_out   (swap_out_0_143),
       .data_out   (data_out_0_143),
       .op_out     (op_out_0_143),
       .pivot_out  (pivot_out_0_143),
       .r          (r_0_143)
     );

  // row 0, col 144

     reg start_in_0_144;
     wire start_out_0_144;

     reg swap_in_0_144;
     wire swap_out_0_144;

     reg [1:0] op_in_0_144;
     wire [1:0] op_out_0_144;

     wire r_0_144;

     wire data_in_0_144;
     wire data_out_0_144;

     reg pivot_in_0_144;
     wire pivot_out_0_144;

     assign data_in_0_144 = data_in[DAT_W-145];

     always @(posedge clk) begin
        op_in_0_144 <= op_out_0_143;
        pivot_in_0_144 <= pivot_out_0_143;
        start_in_0_144 <= start_out_0_143;
        swap_in_0_144 <= swap_out_0_143;
     end
  
     processor_AB AB_0_144 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_144),
       .start_in   (start_in_0_144),
       .swap_in    (swap_in_0_144),
       .op_in      (op_in_0_144),
       .pivot_in   (pivot_in_0_144),
       .start_out  (start_out_0_144),
       .swap_out   (swap_out_0_144),
       .data_out   (data_out_0_144),
       .op_out     (op_out_0_144),
       .pivot_out  (pivot_out_0_144),
       .r          (r_0_144)
     );

  // row 0, col 145

     reg start_in_0_145;
     wire start_out_0_145;

     reg swap_in_0_145;
     wire swap_out_0_145;

     reg [1:0] op_in_0_145;
     wire [1:0] op_out_0_145;

     wire r_0_145;

     wire data_in_0_145;
     wire data_out_0_145;

     reg pivot_in_0_145;
     wire pivot_out_0_145;

     assign data_in_0_145 = data_in[DAT_W-146];

     always @(posedge clk) begin
        op_in_0_145 <= op_out_0_144;
        pivot_in_0_145 <= pivot_out_0_144;
        start_in_0_145 <= start_out_0_144;
        swap_in_0_145 <= swap_out_0_144;
     end
  
     processor_AB AB_0_145 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_145),
       .start_in   (start_in_0_145),
       .swap_in    (swap_in_0_145),
       .op_in      (op_in_0_145),
       .pivot_in   (pivot_in_0_145),
       .start_out  (start_out_0_145),
       .swap_out   (swap_out_0_145),
       .data_out   (data_out_0_145),
       .op_out     (op_out_0_145),
       .pivot_out  (pivot_out_0_145),
       .r          (r_0_145)
     );

  // row 0, col 146

     reg start_in_0_146;
     wire start_out_0_146;

     reg swap_in_0_146;
     wire swap_out_0_146;

     reg [1:0] op_in_0_146;
     wire [1:0] op_out_0_146;

     wire r_0_146;

     wire data_in_0_146;
     wire data_out_0_146;

     reg pivot_in_0_146;
     wire pivot_out_0_146;

     assign data_in_0_146 = data_in[DAT_W-147];

     always @(posedge clk) begin
        op_in_0_146 <= op_out_0_145;
        pivot_in_0_146 <= pivot_out_0_145;
        start_in_0_146 <= start_out_0_145;
        swap_in_0_146 <= swap_out_0_145;
     end
  
     processor_AB AB_0_146 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_146),
       .start_in   (start_in_0_146),
       .swap_in    (swap_in_0_146),
       .op_in      (op_in_0_146),
       .pivot_in   (pivot_in_0_146),
       .start_out  (start_out_0_146),
       .swap_out   (swap_out_0_146),
       .data_out   (data_out_0_146),
       .op_out     (op_out_0_146),
       .pivot_out  (pivot_out_0_146),
       .r          (r_0_146)
     );

  // row 0, col 147

     reg start_in_0_147;
     wire start_out_0_147;

     reg swap_in_0_147;
     wire swap_out_0_147;

     reg [1:0] op_in_0_147;
     wire [1:0] op_out_0_147;

     wire r_0_147;

     wire data_in_0_147;
     wire data_out_0_147;

     reg pivot_in_0_147;
     wire pivot_out_0_147;

     assign data_in_0_147 = data_in[DAT_W-148];

     always @(posedge clk) begin
        op_in_0_147 <= op_out_0_146;
        pivot_in_0_147 <= pivot_out_0_146;
        start_in_0_147 <= start_out_0_146;
        swap_in_0_147 <= swap_out_0_146;
     end
  
     processor_AB AB_0_147 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_147),
       .start_in   (start_in_0_147),
       .swap_in    (swap_in_0_147),
       .op_in      (op_in_0_147),
       .pivot_in   (pivot_in_0_147),
       .start_out  (start_out_0_147),
       .swap_out   (swap_out_0_147),
       .data_out   (data_out_0_147),
       .op_out     (op_out_0_147),
       .pivot_out  (pivot_out_0_147),
       .r          (r_0_147)
     );

  // row 0, col 148

     reg start_in_0_148;
     wire start_out_0_148;

     reg swap_in_0_148;
     wire swap_out_0_148;

     reg [1:0] op_in_0_148;
     wire [1:0] op_out_0_148;

     wire r_0_148;

     wire data_in_0_148;
     wire data_out_0_148;

     reg pivot_in_0_148;
     wire pivot_out_0_148;

     assign data_in_0_148 = data_in[DAT_W-149];

     always @(posedge clk) begin
        op_in_0_148 <= op_out_0_147;
        pivot_in_0_148 <= pivot_out_0_147;
        start_in_0_148 <= start_out_0_147;
        swap_in_0_148 <= swap_out_0_147;
     end
  
     processor_AB AB_0_148 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_148),
       .start_in   (start_in_0_148),
       .swap_in    (swap_in_0_148),
       .op_in      (op_in_0_148),
       .pivot_in   (pivot_in_0_148),
       .start_out  (start_out_0_148),
       .swap_out   (swap_out_0_148),
       .data_out   (data_out_0_148),
       .op_out     (op_out_0_148),
       .pivot_out  (pivot_out_0_148),
       .r          (r_0_148)
     );

  // row 0, col 149

     reg start_in_0_149;
     wire start_out_0_149;

     reg swap_in_0_149;
     wire swap_out_0_149;

     reg [1:0] op_in_0_149;
     wire [1:0] op_out_0_149;

     wire r_0_149;

     wire data_in_0_149;
     wire data_out_0_149;

     reg pivot_in_0_149;
     wire pivot_out_0_149;

     assign data_in_0_149 = data_in[DAT_W-150];

     always @(posedge clk) begin
        op_in_0_149 <= op_out_0_148;
        pivot_in_0_149 <= pivot_out_0_148;
        start_in_0_149 <= start_out_0_148;
        swap_in_0_149 <= swap_out_0_148;
     end
  
     processor_AB AB_0_149 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_149),
       .start_in   (start_in_0_149),
       .swap_in    (swap_in_0_149),
       .op_in      (op_in_0_149),
       .pivot_in   (pivot_in_0_149),
       .start_out  (start_out_0_149),
       .swap_out   (swap_out_0_149),
       .data_out   (data_out_0_149),
       .op_out     (op_out_0_149),
       .pivot_out  (pivot_out_0_149),
       .r          (r_0_149)
     );

  // row 0, col 150

     reg start_in_0_150;
     wire start_out_0_150;

     reg swap_in_0_150;
     wire swap_out_0_150;

     reg [1:0] op_in_0_150;
     wire [1:0] op_out_0_150;

     wire r_0_150;

     wire data_in_0_150;
     wire data_out_0_150;

     reg pivot_in_0_150;
     wire pivot_out_0_150;

     assign data_in_0_150 = data_in[DAT_W-151];

     always @(posedge clk) begin
        op_in_0_150 <= op_out_0_149;
        pivot_in_0_150 <= pivot_out_0_149;
        start_in_0_150 <= start_out_0_149;
        swap_in_0_150 <= swap_out_0_149;
     end
  
     processor_AB AB_0_150 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_150),
       .start_in   (start_in_0_150),
       .swap_in    (swap_in_0_150),
       .op_in      (op_in_0_150),
       .pivot_in   (pivot_in_0_150),
       .start_out  (start_out_0_150),
       .swap_out   (swap_out_0_150),
       .data_out   (data_out_0_150),
       .op_out     (op_out_0_150),
       .pivot_out  (pivot_out_0_150),
       .r          (r_0_150)
     );

  // row 0, col 151

     reg start_in_0_151;
     wire start_out_0_151;

     reg swap_in_0_151;
     wire swap_out_0_151;

     reg [1:0] op_in_0_151;
     wire [1:0] op_out_0_151;

     wire r_0_151;

     wire data_in_0_151;
     wire data_out_0_151;

     reg pivot_in_0_151;
     wire pivot_out_0_151;

     assign data_in_0_151 = data_in[DAT_W-152];

     always @(posedge clk) begin
        op_in_0_151 <= op_out_0_150;
        pivot_in_0_151 <= pivot_out_0_150;
        start_in_0_151 <= start_out_0_150;
        swap_in_0_151 <= swap_out_0_150;
     end
  
     processor_AB AB_0_151 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_151),
       .start_in   (start_in_0_151),
       .swap_in    (swap_in_0_151),
       .op_in      (op_in_0_151),
       .pivot_in   (pivot_in_0_151),
       .start_out  (start_out_0_151),
       .swap_out   (swap_out_0_151),
       .data_out   (data_out_0_151),
       .op_out     (op_out_0_151),
       .pivot_out  (pivot_out_0_151),
       .r          (r_0_151)
     );

  // row 0, col 152

     reg start_in_0_152;
     wire start_out_0_152;

     reg swap_in_0_152;
     wire swap_out_0_152;

     reg [1:0] op_in_0_152;
     wire [1:0] op_out_0_152;

     wire r_0_152;

     wire data_in_0_152;
     wire data_out_0_152;

     reg pivot_in_0_152;
     wire pivot_out_0_152;

     assign data_in_0_152 = data_in[DAT_W-153];

     always @(posedge clk) begin
        op_in_0_152 <= op_out_0_151;
        pivot_in_0_152 <= pivot_out_0_151;
        start_in_0_152 <= start_out_0_151;
        swap_in_0_152 <= swap_out_0_151;
     end
  
     processor_AB AB_0_152 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_152),
       .start_in   (start_in_0_152),
       .swap_in    (swap_in_0_152),
       .op_in      (op_in_0_152),
       .pivot_in   (pivot_in_0_152),
       .start_out  (start_out_0_152),
       .swap_out   (swap_out_0_152),
       .data_out   (data_out_0_152),
       .op_out     (op_out_0_152),
       .pivot_out  (pivot_out_0_152),
       .r          (r_0_152)
     );

  // row 0, col 153

     reg start_in_0_153;
     wire start_out_0_153;

     reg swap_in_0_153;
     wire swap_out_0_153;

     reg [1:0] op_in_0_153;
     wire [1:0] op_out_0_153;

     wire r_0_153;

     wire data_in_0_153;
     wire data_out_0_153;

     reg pivot_in_0_153;
     wire pivot_out_0_153;

     assign data_in_0_153 = data_in[DAT_W-154];

     always @(posedge clk) begin
        op_in_0_153 <= op_out_0_152;
        pivot_in_0_153 <= pivot_out_0_152;
        start_in_0_153 <= start_out_0_152;
        swap_in_0_153 <= swap_out_0_152;
     end
  
     processor_AB AB_0_153 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_153),
       .start_in   (start_in_0_153),
       .swap_in    (swap_in_0_153),
       .op_in      (op_in_0_153),
       .pivot_in   (pivot_in_0_153),
       .start_out  (start_out_0_153),
       .swap_out   (swap_out_0_153),
       .data_out   (data_out_0_153),
       .op_out     (op_out_0_153),
       .pivot_out  (pivot_out_0_153),
       .r          (r_0_153)
     );

  // row 0, col 154

     reg start_in_0_154;
     wire start_out_0_154;

     reg swap_in_0_154;
     wire swap_out_0_154;

     reg [1:0] op_in_0_154;
     wire [1:0] op_out_0_154;

     wire r_0_154;

     wire data_in_0_154;
     wire data_out_0_154;

     reg pivot_in_0_154;
     wire pivot_out_0_154;

     assign data_in_0_154 = data_in[DAT_W-155];

     always @(posedge clk) begin
        op_in_0_154 <= op_out_0_153;
        pivot_in_0_154 <= pivot_out_0_153;
        start_in_0_154 <= start_out_0_153;
        swap_in_0_154 <= swap_out_0_153;
     end
  
     processor_AB AB_0_154 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_154),
       .start_in   (start_in_0_154),
       .swap_in    (swap_in_0_154),
       .op_in      (op_in_0_154),
       .pivot_in   (pivot_in_0_154),
       .start_out  (start_out_0_154),
       .swap_out   (swap_out_0_154),
       .data_out   (data_out_0_154),
       .op_out     (op_out_0_154),
       .pivot_out  (pivot_out_0_154),
       .r          (r_0_154)
     );

  // row 0, col 155

     reg start_in_0_155;
     wire start_out_0_155;

     reg swap_in_0_155;
     wire swap_out_0_155;

     reg [1:0] op_in_0_155;
     wire [1:0] op_out_0_155;

     wire r_0_155;

     wire data_in_0_155;
     wire data_out_0_155;

     reg pivot_in_0_155;
     wire pivot_out_0_155;

     assign data_in_0_155 = data_in[DAT_W-156];

     always @(posedge clk) begin
        op_in_0_155 <= op_out_0_154;
        pivot_in_0_155 <= pivot_out_0_154;
        start_in_0_155 <= start_out_0_154;
        swap_in_0_155 <= swap_out_0_154;
     end
  
     processor_AB AB_0_155 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_155),
       .start_in   (start_in_0_155),
       .swap_in    (swap_in_0_155),
       .op_in      (op_in_0_155),
       .pivot_in   (pivot_in_0_155),
       .start_out  (start_out_0_155),
       .swap_out   (swap_out_0_155),
       .data_out   (data_out_0_155),
       .op_out     (op_out_0_155),
       .pivot_out  (pivot_out_0_155),
       .r          (r_0_155)
     );

  // row 0, col 156

     reg start_in_0_156;
     wire start_out_0_156;

     reg swap_in_0_156;
     wire swap_out_0_156;

     reg [1:0] op_in_0_156;
     wire [1:0] op_out_0_156;

     wire r_0_156;

     wire data_in_0_156;
     wire data_out_0_156;

     reg pivot_in_0_156;
     wire pivot_out_0_156;

     assign data_in_0_156 = data_in[DAT_W-157];

     always @(posedge clk) begin
        op_in_0_156 <= op_out_0_155;
        pivot_in_0_156 <= pivot_out_0_155;
        start_in_0_156 <= start_out_0_155;
        swap_in_0_156 <= swap_out_0_155;
     end
  
     processor_AB AB_0_156 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_156),
       .start_in   (start_in_0_156),
       .swap_in    (swap_in_0_156),
       .op_in      (op_in_0_156),
       .pivot_in   (pivot_in_0_156),
       .start_out  (start_out_0_156),
       .swap_out   (swap_out_0_156),
       .data_out   (data_out_0_156),
       .op_out     (op_out_0_156),
       .pivot_out  (pivot_out_0_156),
       .r          (r_0_156)
     );

  // row 0, col 157

     reg start_in_0_157;
     wire start_out_0_157;

     reg swap_in_0_157;
     wire swap_out_0_157;

     reg [1:0] op_in_0_157;
     wire [1:0] op_out_0_157;

     wire r_0_157;

     wire data_in_0_157;
     wire data_out_0_157;

     reg pivot_in_0_157;
     wire pivot_out_0_157;

     assign data_in_0_157 = data_in[DAT_W-158];

     always @(posedge clk) begin
        op_in_0_157 <= op_out_0_156;
        pivot_in_0_157 <= pivot_out_0_156;
        start_in_0_157 <= start_out_0_156;
        swap_in_0_157 <= swap_out_0_156;
     end
  
     processor_AB AB_0_157 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_157),
       .start_in   (start_in_0_157),
       .swap_in    (swap_in_0_157),
       .op_in      (op_in_0_157),
       .pivot_in   (pivot_in_0_157),
       .start_out  (start_out_0_157),
       .swap_out   (swap_out_0_157),
       .data_out   (data_out_0_157),
       .op_out     (op_out_0_157),
       .pivot_out  (pivot_out_0_157),
       .r          (r_0_157)
     );

  // row 0, col 158

     reg start_in_0_158;
     wire start_out_0_158;

     reg swap_in_0_158;
     wire swap_out_0_158;

     reg [1:0] op_in_0_158;
     wire [1:0] op_out_0_158;

     wire r_0_158;

     wire data_in_0_158;
     wire data_out_0_158;

     reg pivot_in_0_158;
     wire pivot_out_0_158;

     assign data_in_0_158 = data_in[DAT_W-159];

     always @(posedge clk) begin
        op_in_0_158 <= op_out_0_157;
        pivot_in_0_158 <= pivot_out_0_157;
        start_in_0_158 <= start_out_0_157;
        swap_in_0_158 <= swap_out_0_157;
     end
  
     processor_AB AB_0_158 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_158),
       .start_in   (start_in_0_158),
       .swap_in    (swap_in_0_158),
       .op_in      (op_in_0_158),
       .pivot_in   (pivot_in_0_158),
       .start_out  (start_out_0_158),
       .swap_out   (swap_out_0_158),
       .data_out   (data_out_0_158),
       .op_out     (op_out_0_158),
       .pivot_out  (pivot_out_0_158),
       .r          (r_0_158)
     );

  // row 0, col 159

     reg start_in_0_159;
     wire start_out_0_159;

     reg swap_in_0_159;
     wire swap_out_0_159;

     reg [1:0] op_in_0_159;
     wire [1:0] op_out_0_159;

     wire r_0_159;

     wire data_in_0_159;
     wire data_out_0_159;

     reg pivot_in_0_159;
     wire pivot_out_0_159;

     assign data_in_0_159 = data_in[DAT_W-160];

     always @(posedge clk) begin
        op_in_0_159 <= op_out_0_158;
        pivot_in_0_159 <= pivot_out_0_158;
        start_in_0_159 <= start_out_0_158;
        swap_in_0_159 <= swap_out_0_158;
     end
  
     processor_AB AB_0_159 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_159),
       .start_in   (start_in_0_159),
       .swap_in    (swap_in_0_159),
       .op_in      (op_in_0_159),
       .pivot_in   (pivot_in_0_159),
       .start_out  (start_out_0_159),
       .swap_out   (swap_out_0_159),
       .data_out   (data_out_0_159),
       .op_out     (op_out_0_159),
       .pivot_out  (pivot_out_0_159),
       .r          (r_0_159)
     );

  // row 0, col 160

     reg start_in_0_160;
     wire start_out_0_160;

     reg swap_in_0_160;
     wire swap_out_0_160;

     reg [1:0] op_in_0_160;
     wire [1:0] op_out_0_160;

     wire r_0_160;

     wire data_in_0_160;
     wire data_out_0_160;

     reg pivot_in_0_160;
     wire pivot_out_0_160;

     assign data_in_0_160 = data_in[DAT_W-161];

     always @(posedge clk) begin
        op_in_0_160 <= op_out_0_159;
        pivot_in_0_160 <= pivot_out_0_159;
        start_in_0_160 <= start_out_0_159;
        swap_in_0_160 <= swap_out_0_159;
     end
  
     processor_AB AB_0_160 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_160),
       .start_in   (start_in_0_160),
       .swap_in    (swap_in_0_160),
       .op_in      (op_in_0_160),
       .pivot_in   (pivot_in_0_160),
       .start_out  (start_out_0_160),
       .swap_out   (swap_out_0_160),
       .data_out   (data_out_0_160),
       .op_out     (op_out_0_160),
       .pivot_out  (pivot_out_0_160),
       .r          (r_0_160)
     );

  // row 0, col 161

     reg start_in_0_161;
     wire start_out_0_161;

     reg swap_in_0_161;
     wire swap_out_0_161;

     reg [1:0] op_in_0_161;
     wire [1:0] op_out_0_161;

     wire r_0_161;

     wire data_in_0_161;
     wire data_out_0_161;

     reg pivot_in_0_161;
     wire pivot_out_0_161;

     assign data_in_0_161 = data_in[DAT_W-162];

     always @(posedge clk) begin
        op_in_0_161 <= op_out_0_160;
        pivot_in_0_161 <= pivot_out_0_160;
        start_in_0_161 <= start_out_0_160;
        swap_in_0_161 <= swap_out_0_160;
     end
  
     processor_AB AB_0_161 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_161),
       .start_in   (start_in_0_161),
       .swap_in    (swap_in_0_161),
       .op_in      (op_in_0_161),
       .pivot_in   (pivot_in_0_161),
       .start_out  (start_out_0_161),
       .swap_out   (swap_out_0_161),
       .data_out   (data_out_0_161),
       .op_out     (op_out_0_161),
       .pivot_out  (pivot_out_0_161),
       .r          (r_0_161)
     );

  // row 0, col 162

     reg start_in_0_162;
     wire start_out_0_162;

     reg swap_in_0_162;
     wire swap_out_0_162;

     reg [1:0] op_in_0_162;
     wire [1:0] op_out_0_162;

     wire r_0_162;

     wire data_in_0_162;
     wire data_out_0_162;

     reg pivot_in_0_162;
     wire pivot_out_0_162;

     assign data_in_0_162 = data_in[DAT_W-163];

     always @(posedge clk) begin
        op_in_0_162 <= op_out_0_161;
        pivot_in_0_162 <= pivot_out_0_161;
        start_in_0_162 <= start_out_0_161;
        swap_in_0_162 <= swap_out_0_161;
     end
  
     processor_AB AB_0_162 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_162),
       .start_in   (start_in_0_162),
       .swap_in    (swap_in_0_162),
       .op_in      (op_in_0_162),
       .pivot_in   (pivot_in_0_162),
       .start_out  (start_out_0_162),
       .swap_out   (swap_out_0_162),
       .data_out   (data_out_0_162),
       .op_out     (op_out_0_162),
       .pivot_out  (pivot_out_0_162),
       .r          (r_0_162)
     );

  // row 0, col 163

     reg start_in_0_163;
     wire start_out_0_163;

     reg swap_in_0_163;
     wire swap_out_0_163;

     reg [1:0] op_in_0_163;
     wire [1:0] op_out_0_163;

     wire r_0_163;

     wire data_in_0_163;
     wire data_out_0_163;

     reg pivot_in_0_163;
     wire pivot_out_0_163;

     assign data_in_0_163 = data_in[DAT_W-164];

     always @(posedge clk) begin
        op_in_0_163 <= op_out_0_162;
        pivot_in_0_163 <= pivot_out_0_162;
        start_in_0_163 <= start_out_0_162;
        swap_in_0_163 <= swap_out_0_162;
     end
  
     processor_AB AB_0_163 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_163),
       .start_in   (start_in_0_163),
       .swap_in    (swap_in_0_163),
       .op_in      (op_in_0_163),
       .pivot_in   (pivot_in_0_163),
       .start_out  (start_out_0_163),
       .swap_out   (swap_out_0_163),
       .data_out   (data_out_0_163),
       .op_out     (op_out_0_163),
       .pivot_out  (pivot_out_0_163),
       .r          (r_0_163)
     );

  // row 0, col 164

     reg start_in_0_164;
     wire start_out_0_164;

     reg swap_in_0_164;
     wire swap_out_0_164;

     reg [1:0] op_in_0_164;
     wire [1:0] op_out_0_164;

     wire r_0_164;

     wire data_in_0_164;
     wire data_out_0_164;

     reg pivot_in_0_164;
     wire pivot_out_0_164;

     assign data_in_0_164 = data_in[DAT_W-165];

     always @(posedge clk) begin
        op_in_0_164 <= op_out_0_163;
        pivot_in_0_164 <= pivot_out_0_163;
        start_in_0_164 <= start_out_0_163;
        swap_in_0_164 <= swap_out_0_163;
     end
  
     processor_AB AB_0_164 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_164),
       .start_in   (start_in_0_164),
       .swap_in    (swap_in_0_164),
       .op_in      (op_in_0_164),
       .pivot_in   (pivot_in_0_164),
       .start_out  (start_out_0_164),
       .swap_out   (swap_out_0_164),
       .data_out   (data_out_0_164),
       .op_out     (op_out_0_164),
       .pivot_out  (pivot_out_0_164),
       .r          (r_0_164)
     );

  // row 0, col 165

     reg start_in_0_165;
     wire start_out_0_165;

     reg swap_in_0_165;
     wire swap_out_0_165;

     reg [1:0] op_in_0_165;
     wire [1:0] op_out_0_165;

     wire r_0_165;

     wire data_in_0_165;
     wire data_out_0_165;

     reg pivot_in_0_165;
     wire pivot_out_0_165;

     assign data_in_0_165 = data_in[DAT_W-166];

     always @(posedge clk) begin
        op_in_0_165 <= op_out_0_164;
        pivot_in_0_165 <= pivot_out_0_164;
        start_in_0_165 <= start_out_0_164;
        swap_in_0_165 <= swap_out_0_164;
     end
  
     processor_AB AB_0_165 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_0_165),
       .start_in   (start_in_0_165),
       .swap_in    (swap_in_0_165),
       .op_in      (op_in_0_165),
       .pivot_in   (pivot_in_0_165),
       .start_out  (start_out_0_165),
       .swap_out   (swap_out_0_165),
       .data_out   (data_out_0_165),
       .op_out     (op_out_0_165),
       .pivot_out  (pivot_out_0_165),
       .r          (r_0_165)
     );

  /////////////////////////////////////
  // row 1
  // row 1, col 0

     wire start_in_1_0;
     wire start_out_1_0;

     wire swap_in_1_0;
     wire swap_out_1_0;

     wire [1:0] op_in_1_0;
     wire [1:0] op_out_1_0;

     wire r_1_0;

     reg data_in_1_0;
     wire data_out_1_0;

     wire pivot_in_1_0;
     wire pivout_out_1_0;

     assign op_in_1_0 = 2'b00;
     assign pivot_in_1_0 = 0;

     assign start_in_1_0 = start_row[1]; 
     assign swap_in_1_0 = mode ? swap : swap_row[1]; 

     always @(posedge clk) begin
         data_in_1_0 <= data_out_0_0;
     end

     processor_AB AB_1_0 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_0),
       .start_in   (start_in_1_0),
       .swap_in   (swap_in_1_0),
       .op_in      (op_in_1_0),
       .pivot_in   (pivot_in_1_0),
       .start_out  (start_out_1_0),
       .swap_out   (swap_out_1_0),
       .data_out   (data_out_1_0),
       .op_out     (op_out_1_0),
       .pivot_out  (pivot_out_1_0),
       .r          (r_1_0)
     );

  // row 1, col 1

     reg start_in_1_1;
     wire start_out_1_1;

     reg swap_in_1_1;
     wire swap_out_1_1;

     reg [1:0] op_in_1_1;
     wire [1:0] op_out_1_1;

     wire r_1_1;

     reg data_in_1_1;
     wire data_out_1_1;

     reg pivot_in_1_1;
     wire pivot_out_1_1;

     always @(posedge clk) begin
         op_in_1_1 <= op_out_1_0;
         pivot_in_1_1 <= pivot_out_1_0;
         start_in_1_1 <= start_out_1_0;
         swap_in_1_1 <= swap_out_1_0;
     end

     always @(posedge clk) begin
         data_in_1_1 <= data_out_0_1;
     end
  
     processor_AB AB_1_1 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_1),
       .start_in   (start_in_1_1),
       .swap_in   (swap_in_1_1),
       .op_in      (op_in_1_1),
       .pivot_in   (pivot_in_1_1),
       .start_out  (start_out_1_1),
       .swap_out   (swap_out_1_1),
       .data_out   (data_out_1_1),
       .op_out     (op_out_1_1),
       .pivot_out  (pivot_out_1_1),
       .r          (r_1_1)
     );

  // row 1, col 2

     reg start_in_1_2;
     wire start_out_1_2;

     reg swap_in_1_2;
     wire swap_out_1_2;

     reg [1:0] op_in_1_2;
     wire [1:0] op_out_1_2;

     wire r_1_2;

     reg data_in_1_2;
     wire data_out_1_2;

     reg pivot_in_1_2;
     wire pivot_out_1_2;

     always @(posedge clk) begin
         op_in_1_2 <= op_out_1_1;
         pivot_in_1_2 <= pivot_out_1_1;
         start_in_1_2 <= start_out_1_1;
         swap_in_1_2 <= swap_out_1_1;
     end

     always @(posedge clk) begin
         data_in_1_2 <= data_out_0_2;
     end
  
     processor_AB AB_1_2 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_2),
       .start_in   (start_in_1_2),
       .swap_in   (swap_in_1_2),
       .op_in      (op_in_1_2),
       .pivot_in   (pivot_in_1_2),
       .start_out  (start_out_1_2),
       .swap_out   (swap_out_1_2),
       .data_out   (data_out_1_2),
       .op_out     (op_out_1_2),
       .pivot_out  (pivot_out_1_2),
       .r          (r_1_2)
     );

  // row 1, col 3

     reg start_in_1_3;
     wire start_out_1_3;

     reg swap_in_1_3;
     wire swap_out_1_3;

     reg [1:0] op_in_1_3;
     wire [1:0] op_out_1_3;

     wire r_1_3;

     reg data_in_1_3;
     wire data_out_1_3;

     reg pivot_in_1_3;
     wire pivot_out_1_3;

     always @(posedge clk) begin
         op_in_1_3 <= op_out_1_2;
         pivot_in_1_3 <= pivot_out_1_2;
         start_in_1_3 <= start_out_1_2;
         swap_in_1_3 <= swap_out_1_2;
     end

     always @(posedge clk) begin
         data_in_1_3 <= data_out_0_3;
     end
  
     processor_AB AB_1_3 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_3),
       .start_in   (start_in_1_3),
       .swap_in   (swap_in_1_3),
       .op_in      (op_in_1_3),
       .pivot_in   (pivot_in_1_3),
       .start_out  (start_out_1_3),
       .swap_out   (swap_out_1_3),
       .data_out   (data_out_1_3),
       .op_out     (op_out_1_3),
       .pivot_out  (pivot_out_1_3),
       .r          (r_1_3)
     );

  // row 1, col 4

     reg start_in_1_4;
     wire start_out_1_4;

     reg swap_in_1_4;
     wire swap_out_1_4;

     reg [1:0] op_in_1_4;
     wire [1:0] op_out_1_4;

     wire r_1_4;

     reg data_in_1_4;
     wire data_out_1_4;

     reg pivot_in_1_4;
     wire pivot_out_1_4;

     always @(posedge clk) begin
         op_in_1_4 <= op_out_1_3;
         pivot_in_1_4 <= pivot_out_1_3;
         start_in_1_4 <= start_out_1_3;
         swap_in_1_4 <= swap_out_1_3;
     end

     always @(posedge clk) begin
         data_in_1_4 <= data_out_0_4;
     end
  
     processor_AB AB_1_4 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_4),
       .start_in   (start_in_1_4),
       .swap_in   (swap_in_1_4),
       .op_in      (op_in_1_4),
       .pivot_in   (pivot_in_1_4),
       .start_out  (start_out_1_4),
       .swap_out   (swap_out_1_4),
       .data_out   (data_out_1_4),
       .op_out     (op_out_1_4),
       .pivot_out  (pivot_out_1_4),
       .r          (r_1_4)
     );

  // row 1, col 5

     reg start_in_1_5;
     wire start_out_1_5;

     reg swap_in_1_5;
     wire swap_out_1_5;

     reg [1:0] op_in_1_5;
     wire [1:0] op_out_1_5;

     wire r_1_5;

     reg data_in_1_5;
     wire data_out_1_5;

     reg pivot_in_1_5;
     wire pivot_out_1_5;

     always @(posedge clk) begin
         op_in_1_5 <= op_out_1_4;
         pivot_in_1_5 <= pivot_out_1_4;
         start_in_1_5 <= start_out_1_4;
         swap_in_1_5 <= swap_out_1_4;
     end

     always @(posedge clk) begin
         data_in_1_5 <= data_out_0_5;
     end
  
     processor_AB AB_1_5 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_5),
       .start_in   (start_in_1_5),
       .swap_in   (swap_in_1_5),
       .op_in      (op_in_1_5),
       .pivot_in   (pivot_in_1_5),
       .start_out  (start_out_1_5),
       .swap_out   (swap_out_1_5),
       .data_out   (data_out_1_5),
       .op_out     (op_out_1_5),
       .pivot_out  (pivot_out_1_5),
       .r          (r_1_5)
     );

  // row 1, col 6

     reg start_in_1_6;
     wire start_out_1_6;

     reg swap_in_1_6;
     wire swap_out_1_6;

     reg [1:0] op_in_1_6;
     wire [1:0] op_out_1_6;

     wire r_1_6;

     reg data_in_1_6;
     wire data_out_1_6;

     reg pivot_in_1_6;
     wire pivot_out_1_6;

     always @(posedge clk) begin
         op_in_1_6 <= op_out_1_5;
         pivot_in_1_6 <= pivot_out_1_5;
         start_in_1_6 <= start_out_1_5;
         swap_in_1_6 <= swap_out_1_5;
     end

     always @(posedge clk) begin
         data_in_1_6 <= data_out_0_6;
     end
  
     processor_AB AB_1_6 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_6),
       .start_in   (start_in_1_6),
       .swap_in   (swap_in_1_6),
       .op_in      (op_in_1_6),
       .pivot_in   (pivot_in_1_6),
       .start_out  (start_out_1_6),
       .swap_out   (swap_out_1_6),
       .data_out   (data_out_1_6),
       .op_out     (op_out_1_6),
       .pivot_out  (pivot_out_1_6),
       .r          (r_1_6)
     );

  // row 1, col 7

     reg start_in_1_7;
     wire start_out_1_7;

     reg swap_in_1_7;
     wire swap_out_1_7;

     reg [1:0] op_in_1_7;
     wire [1:0] op_out_1_7;

     wire r_1_7;

     reg data_in_1_7;
     wire data_out_1_7;

     reg pivot_in_1_7;
     wire pivot_out_1_7;

     always @(posedge clk) begin
         op_in_1_7 <= op_out_1_6;
         pivot_in_1_7 <= pivot_out_1_6;
         start_in_1_7 <= start_out_1_6;
         swap_in_1_7 <= swap_out_1_6;
     end

     always @(posedge clk) begin
         data_in_1_7 <= data_out_0_7;
     end
  
     processor_AB AB_1_7 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_7),
       .start_in   (start_in_1_7),
       .swap_in   (swap_in_1_7),
       .op_in      (op_in_1_7),
       .pivot_in   (pivot_in_1_7),
       .start_out  (start_out_1_7),
       .swap_out   (swap_out_1_7),
       .data_out   (data_out_1_7),
       .op_out     (op_out_1_7),
       .pivot_out  (pivot_out_1_7),
       .r          (r_1_7)
     );

  // row 1, col 8

     reg start_in_1_8;
     wire start_out_1_8;

     reg swap_in_1_8;
     wire swap_out_1_8;

     reg [1:0] op_in_1_8;
     wire [1:0] op_out_1_8;

     wire r_1_8;

     reg data_in_1_8;
     wire data_out_1_8;

     reg pivot_in_1_8;
     wire pivot_out_1_8;

     always @(posedge clk) begin
         op_in_1_8 <= op_out_1_7;
         pivot_in_1_8 <= pivot_out_1_7;
         start_in_1_8 <= start_out_1_7;
         swap_in_1_8 <= swap_out_1_7;
     end

     always @(posedge clk) begin
         data_in_1_8 <= data_out_0_8;
     end
  
     processor_AB AB_1_8 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_8),
       .start_in   (start_in_1_8),
       .swap_in   (swap_in_1_8),
       .op_in      (op_in_1_8),
       .pivot_in   (pivot_in_1_8),
       .start_out  (start_out_1_8),
       .swap_out   (swap_out_1_8),
       .data_out   (data_out_1_8),
       .op_out     (op_out_1_8),
       .pivot_out  (pivot_out_1_8),
       .r          (r_1_8)
     );

  // row 1, col 9

     reg start_in_1_9;
     wire start_out_1_9;

     reg swap_in_1_9;
     wire swap_out_1_9;

     reg [1:0] op_in_1_9;
     wire [1:0] op_out_1_9;

     wire r_1_9;

     reg data_in_1_9;
     wire data_out_1_9;

     reg pivot_in_1_9;
     wire pivot_out_1_9;

     always @(posedge clk) begin
         op_in_1_9 <= op_out_1_8;
         pivot_in_1_9 <= pivot_out_1_8;
         start_in_1_9 <= start_out_1_8;
         swap_in_1_9 <= swap_out_1_8;
     end

     always @(posedge clk) begin
         data_in_1_9 <= data_out_0_9;
     end
  
     processor_AB AB_1_9 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_9),
       .start_in   (start_in_1_9),
       .swap_in   (swap_in_1_9),
       .op_in      (op_in_1_9),
       .pivot_in   (pivot_in_1_9),
       .start_out  (start_out_1_9),
       .swap_out   (swap_out_1_9),
       .data_out   (data_out_1_9),
       .op_out     (op_out_1_9),
       .pivot_out  (pivot_out_1_9),
       .r          (r_1_9)
     );

  // row 1, col 10

     reg start_in_1_10;
     wire start_out_1_10;

     reg swap_in_1_10;
     wire swap_out_1_10;

     reg [1:0] op_in_1_10;
     wire [1:0] op_out_1_10;

     wire r_1_10;

     reg data_in_1_10;
     wire data_out_1_10;

     reg pivot_in_1_10;
     wire pivot_out_1_10;

     always @(posedge clk) begin
         op_in_1_10 <= op_out_1_9;
         pivot_in_1_10 <= pivot_out_1_9;
         start_in_1_10 <= start_out_1_9;
         swap_in_1_10 <= swap_out_1_9;
     end

     always @(posedge clk) begin
         data_in_1_10 <= data_out_0_10;
     end
  
     processor_AB AB_1_10 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_10),
       .start_in   (start_in_1_10),
       .swap_in   (swap_in_1_10),
       .op_in      (op_in_1_10),
       .pivot_in   (pivot_in_1_10),
       .start_out  (start_out_1_10),
       .swap_out   (swap_out_1_10),
       .data_out   (data_out_1_10),
       .op_out     (op_out_1_10),
       .pivot_out  (pivot_out_1_10),
       .r          (r_1_10)
     );

  // row 1, col 11

     reg start_in_1_11;
     wire start_out_1_11;

     reg swap_in_1_11;
     wire swap_out_1_11;

     reg [1:0] op_in_1_11;
     wire [1:0] op_out_1_11;

     wire r_1_11;

     reg data_in_1_11;
     wire data_out_1_11;

     reg pivot_in_1_11;
     wire pivot_out_1_11;

     always @(posedge clk) begin
         op_in_1_11 <= op_out_1_10;
         pivot_in_1_11 <= pivot_out_1_10;
         start_in_1_11 <= start_out_1_10;
         swap_in_1_11 <= swap_out_1_10;
     end

     always @(posedge clk) begin
         data_in_1_11 <= data_out_0_11;
     end
  
     processor_AB AB_1_11 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_11),
       .start_in   (start_in_1_11),
       .swap_in   (swap_in_1_11),
       .op_in      (op_in_1_11),
       .pivot_in   (pivot_in_1_11),
       .start_out  (start_out_1_11),
       .swap_out   (swap_out_1_11),
       .data_out   (data_out_1_11),
       .op_out     (op_out_1_11),
       .pivot_out  (pivot_out_1_11),
       .r          (r_1_11)
     );

  // row 1, col 12

     reg start_in_1_12;
     wire start_out_1_12;

     reg swap_in_1_12;
     wire swap_out_1_12;

     reg [1:0] op_in_1_12;
     wire [1:0] op_out_1_12;

     wire r_1_12;

     reg data_in_1_12;
     wire data_out_1_12;

     reg pivot_in_1_12;
     wire pivot_out_1_12;

     always @(posedge clk) begin
         op_in_1_12 <= op_out_1_11;
         pivot_in_1_12 <= pivot_out_1_11;
         start_in_1_12 <= start_out_1_11;
         swap_in_1_12 <= swap_out_1_11;
     end

     always @(posedge clk) begin
         data_in_1_12 <= data_out_0_12;
     end
  
     processor_AB AB_1_12 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_12),
       .start_in   (start_in_1_12),
       .swap_in   (swap_in_1_12),
       .op_in      (op_in_1_12),
       .pivot_in   (pivot_in_1_12),
       .start_out  (start_out_1_12),
       .swap_out   (swap_out_1_12),
       .data_out   (data_out_1_12),
       .op_out     (op_out_1_12),
       .pivot_out  (pivot_out_1_12),
       .r          (r_1_12)
     );

  // row 1, col 13

     reg start_in_1_13;
     wire start_out_1_13;

     reg swap_in_1_13;
     wire swap_out_1_13;

     reg [1:0] op_in_1_13;
     wire [1:0] op_out_1_13;

     wire r_1_13;

     reg data_in_1_13;
     wire data_out_1_13;

     reg pivot_in_1_13;
     wire pivot_out_1_13;

     always @(posedge clk) begin
         op_in_1_13 <= op_out_1_12;
         pivot_in_1_13 <= pivot_out_1_12;
         start_in_1_13 <= start_out_1_12;
         swap_in_1_13 <= swap_out_1_12;
     end

     always @(posedge clk) begin
         data_in_1_13 <= data_out_0_13;
     end
  
     processor_AB AB_1_13 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_13),
       .start_in   (start_in_1_13),
       .swap_in   (swap_in_1_13),
       .op_in      (op_in_1_13),
       .pivot_in   (pivot_in_1_13),
       .start_out  (start_out_1_13),
       .swap_out   (swap_out_1_13),
       .data_out   (data_out_1_13),
       .op_out     (op_out_1_13),
       .pivot_out  (pivot_out_1_13),
       .r          (r_1_13)
     );

  // row 1, col 14

     reg start_in_1_14;
     wire start_out_1_14;

     reg swap_in_1_14;
     wire swap_out_1_14;

     reg [1:0] op_in_1_14;
     wire [1:0] op_out_1_14;

     wire r_1_14;

     reg data_in_1_14;
     wire data_out_1_14;

     reg pivot_in_1_14;
     wire pivot_out_1_14;

     always @(posedge clk) begin
         op_in_1_14 <= op_out_1_13;
         pivot_in_1_14 <= pivot_out_1_13;
         start_in_1_14 <= start_out_1_13;
         swap_in_1_14 <= swap_out_1_13;
     end

     always @(posedge clk) begin
         data_in_1_14 <= data_out_0_14;
     end
  
     processor_AB AB_1_14 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_14),
       .start_in   (start_in_1_14),
       .swap_in   (swap_in_1_14),
       .op_in      (op_in_1_14),
       .pivot_in   (pivot_in_1_14),
       .start_out  (start_out_1_14),
       .swap_out   (swap_out_1_14),
       .data_out   (data_out_1_14),
       .op_out     (op_out_1_14),
       .pivot_out  (pivot_out_1_14),
       .r          (r_1_14)
     );

  // row 1, col 15

     reg start_in_1_15;
     wire start_out_1_15;

     reg swap_in_1_15;
     wire swap_out_1_15;

     reg [1:0] op_in_1_15;
     wire [1:0] op_out_1_15;

     wire r_1_15;

     reg data_in_1_15;
     wire data_out_1_15;

     reg pivot_in_1_15;
     wire pivot_out_1_15;

     always @(posedge clk) begin
         op_in_1_15 <= op_out_1_14;
         pivot_in_1_15 <= pivot_out_1_14;
         start_in_1_15 <= start_out_1_14;
         swap_in_1_15 <= swap_out_1_14;
     end

     always @(posedge clk) begin
         data_in_1_15 <= data_out_0_15;
     end
  
     processor_AB AB_1_15 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_15),
       .start_in   (start_in_1_15),
       .swap_in   (swap_in_1_15),
       .op_in      (op_in_1_15),
       .pivot_in   (pivot_in_1_15),
       .start_out  (start_out_1_15),
       .swap_out   (swap_out_1_15),
       .data_out   (data_out_1_15),
       .op_out     (op_out_1_15),
       .pivot_out  (pivot_out_1_15),
       .r          (r_1_15)
     );

  // row 1, col 16

     reg start_in_1_16;
     wire start_out_1_16;

     reg swap_in_1_16;
     wire swap_out_1_16;

     reg [1:0] op_in_1_16;
     wire [1:0] op_out_1_16;

     wire r_1_16;

     reg data_in_1_16;
     wire data_out_1_16;

     reg pivot_in_1_16;
     wire pivot_out_1_16;

     always @(posedge clk) begin
         op_in_1_16 <= op_out_1_15;
         pivot_in_1_16 <= pivot_out_1_15;
         start_in_1_16 <= start_out_1_15;
         swap_in_1_16 <= swap_out_1_15;
     end

     always @(posedge clk) begin
         data_in_1_16 <= data_out_0_16;
     end
  
     processor_AB AB_1_16 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_16),
       .start_in   (start_in_1_16),
       .swap_in   (swap_in_1_16),
       .op_in      (op_in_1_16),
       .pivot_in   (pivot_in_1_16),
       .start_out  (start_out_1_16),
       .swap_out   (swap_out_1_16),
       .data_out   (data_out_1_16),
       .op_out     (op_out_1_16),
       .pivot_out  (pivot_out_1_16),
       .r          (r_1_16)
     );

  // row 1, col 17

     reg start_in_1_17;
     wire start_out_1_17;

     reg swap_in_1_17;
     wire swap_out_1_17;

     reg [1:0] op_in_1_17;
     wire [1:0] op_out_1_17;

     wire r_1_17;

     reg data_in_1_17;
     wire data_out_1_17;

     reg pivot_in_1_17;
     wire pivot_out_1_17;

     always @(posedge clk) begin
         op_in_1_17 <= op_out_1_16;
         pivot_in_1_17 <= pivot_out_1_16;
         start_in_1_17 <= start_out_1_16;
         swap_in_1_17 <= swap_out_1_16;
     end

     always @(posedge clk) begin
         data_in_1_17 <= data_out_0_17;
     end
  
     processor_AB AB_1_17 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_17),
       .start_in   (start_in_1_17),
       .swap_in   (swap_in_1_17),
       .op_in      (op_in_1_17),
       .pivot_in   (pivot_in_1_17),
       .start_out  (start_out_1_17),
       .swap_out   (swap_out_1_17),
       .data_out   (data_out_1_17),
       .op_out     (op_out_1_17),
       .pivot_out  (pivot_out_1_17),
       .r          (r_1_17)
     );

  // row 1, col 18

     reg start_in_1_18;
     wire start_out_1_18;

     reg swap_in_1_18;
     wire swap_out_1_18;

     reg [1:0] op_in_1_18;
     wire [1:0] op_out_1_18;

     wire r_1_18;

     reg data_in_1_18;
     wire data_out_1_18;

     reg pivot_in_1_18;
     wire pivot_out_1_18;

     always @(posedge clk) begin
         op_in_1_18 <= op_out_1_17;
         pivot_in_1_18 <= pivot_out_1_17;
         start_in_1_18 <= start_out_1_17;
         swap_in_1_18 <= swap_out_1_17;
     end

     always @(posedge clk) begin
         data_in_1_18 <= data_out_0_18;
     end
  
     processor_AB AB_1_18 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_18),
       .start_in   (start_in_1_18),
       .swap_in   (swap_in_1_18),
       .op_in      (op_in_1_18),
       .pivot_in   (pivot_in_1_18),
       .start_out  (start_out_1_18),
       .swap_out   (swap_out_1_18),
       .data_out   (data_out_1_18),
       .op_out     (op_out_1_18),
       .pivot_out  (pivot_out_1_18),
       .r          (r_1_18)
     );

  // row 1, col 19

     reg start_in_1_19;
     wire start_out_1_19;

     reg swap_in_1_19;
     wire swap_out_1_19;

     reg [1:0] op_in_1_19;
     wire [1:0] op_out_1_19;

     wire r_1_19;

     reg data_in_1_19;
     wire data_out_1_19;

     reg pivot_in_1_19;
     wire pivot_out_1_19;

     always @(posedge clk) begin
         op_in_1_19 <= op_out_1_18;
         pivot_in_1_19 <= pivot_out_1_18;
         start_in_1_19 <= start_out_1_18;
         swap_in_1_19 <= swap_out_1_18;
     end

     always @(posedge clk) begin
         data_in_1_19 <= data_out_0_19;
     end
  
     processor_AB AB_1_19 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_19),
       .start_in   (start_in_1_19),
       .swap_in   (swap_in_1_19),
       .op_in      (op_in_1_19),
       .pivot_in   (pivot_in_1_19),
       .start_out  (start_out_1_19),
       .swap_out   (swap_out_1_19),
       .data_out   (data_out_1_19),
       .op_out     (op_out_1_19),
       .pivot_out  (pivot_out_1_19),
       .r          (r_1_19)
     );

  // row 1, col 20

     reg start_in_1_20;
     wire start_out_1_20;

     reg swap_in_1_20;
     wire swap_out_1_20;

     reg [1:0] op_in_1_20;
     wire [1:0] op_out_1_20;

     wire r_1_20;

     reg data_in_1_20;
     wire data_out_1_20;

     reg pivot_in_1_20;
     wire pivot_out_1_20;

     always @(posedge clk) begin
         op_in_1_20 <= op_out_1_19;
         pivot_in_1_20 <= pivot_out_1_19;
         start_in_1_20 <= start_out_1_19;
         swap_in_1_20 <= swap_out_1_19;
     end

     always @(posedge clk) begin
         data_in_1_20 <= data_out_0_20;
     end
  
     processor_AB AB_1_20 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_20),
       .start_in   (start_in_1_20),
       .swap_in   (swap_in_1_20),
       .op_in      (op_in_1_20),
       .pivot_in   (pivot_in_1_20),
       .start_out  (start_out_1_20),
       .swap_out   (swap_out_1_20),
       .data_out   (data_out_1_20),
       .op_out     (op_out_1_20),
       .pivot_out  (pivot_out_1_20),
       .r          (r_1_20)
     );

  // row 1, col 21

     reg start_in_1_21;
     wire start_out_1_21;

     reg swap_in_1_21;
     wire swap_out_1_21;

     reg [1:0] op_in_1_21;
     wire [1:0] op_out_1_21;

     wire r_1_21;

     reg data_in_1_21;
     wire data_out_1_21;

     reg pivot_in_1_21;
     wire pivot_out_1_21;

     always @(posedge clk) begin
         op_in_1_21 <= op_out_1_20;
         pivot_in_1_21 <= pivot_out_1_20;
         start_in_1_21 <= start_out_1_20;
         swap_in_1_21 <= swap_out_1_20;
     end

     always @(posedge clk) begin
         data_in_1_21 <= data_out_0_21;
     end
  
     processor_AB AB_1_21 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_21),
       .start_in   (start_in_1_21),
       .swap_in   (swap_in_1_21),
       .op_in      (op_in_1_21),
       .pivot_in   (pivot_in_1_21),
       .start_out  (start_out_1_21),
       .swap_out   (swap_out_1_21),
       .data_out   (data_out_1_21),
       .op_out     (op_out_1_21),
       .pivot_out  (pivot_out_1_21),
       .r          (r_1_21)
     );

  // row 1, col 22

     reg start_in_1_22;
     wire start_out_1_22;

     reg swap_in_1_22;
     wire swap_out_1_22;

     reg [1:0] op_in_1_22;
     wire [1:0] op_out_1_22;

     wire r_1_22;

     reg data_in_1_22;
     wire data_out_1_22;

     reg pivot_in_1_22;
     wire pivot_out_1_22;

     always @(posedge clk) begin
         op_in_1_22 <= op_out_1_21;
         pivot_in_1_22 <= pivot_out_1_21;
         start_in_1_22 <= start_out_1_21;
         swap_in_1_22 <= swap_out_1_21;
     end

     always @(posedge clk) begin
         data_in_1_22 <= data_out_0_22;
     end
  
     processor_AB AB_1_22 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_22),
       .start_in   (start_in_1_22),
       .swap_in   (swap_in_1_22),
       .op_in      (op_in_1_22),
       .pivot_in   (pivot_in_1_22),
       .start_out  (start_out_1_22),
       .swap_out   (swap_out_1_22),
       .data_out   (data_out_1_22),
       .op_out     (op_out_1_22),
       .pivot_out  (pivot_out_1_22),
       .r          (r_1_22)
     );

  // row 1, col 23

     reg start_in_1_23;
     wire start_out_1_23;

     reg swap_in_1_23;
     wire swap_out_1_23;

     reg [1:0] op_in_1_23;
     wire [1:0] op_out_1_23;

     wire r_1_23;

     reg data_in_1_23;
     wire data_out_1_23;

     reg pivot_in_1_23;
     wire pivot_out_1_23;

     always @(posedge clk) begin
         op_in_1_23 <= op_out_1_22;
         pivot_in_1_23 <= pivot_out_1_22;
         start_in_1_23 <= start_out_1_22;
         swap_in_1_23 <= swap_out_1_22;
     end

     always @(posedge clk) begin
         data_in_1_23 <= data_out_0_23;
     end
  
     processor_AB AB_1_23 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_23),
       .start_in   (start_in_1_23),
       .swap_in   (swap_in_1_23),
       .op_in      (op_in_1_23),
       .pivot_in   (pivot_in_1_23),
       .start_out  (start_out_1_23),
       .swap_out   (swap_out_1_23),
       .data_out   (data_out_1_23),
       .op_out     (op_out_1_23),
       .pivot_out  (pivot_out_1_23),
       .r          (r_1_23)
     );

  // row 1, col 24

     reg start_in_1_24;
     wire start_out_1_24;

     reg swap_in_1_24;
     wire swap_out_1_24;

     reg [1:0] op_in_1_24;
     wire [1:0] op_out_1_24;

     wire r_1_24;

     reg data_in_1_24;
     wire data_out_1_24;

     reg pivot_in_1_24;
     wire pivot_out_1_24;

     always @(posedge clk) begin
         op_in_1_24 <= op_out_1_23;
         pivot_in_1_24 <= pivot_out_1_23;
         start_in_1_24 <= start_out_1_23;
         swap_in_1_24 <= swap_out_1_23;
     end

     always @(posedge clk) begin
         data_in_1_24 <= data_out_0_24;
     end
  
     processor_AB AB_1_24 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_24),
       .start_in   (start_in_1_24),
       .swap_in   (swap_in_1_24),
       .op_in      (op_in_1_24),
       .pivot_in   (pivot_in_1_24),
       .start_out  (start_out_1_24),
       .swap_out   (swap_out_1_24),
       .data_out   (data_out_1_24),
       .op_out     (op_out_1_24),
       .pivot_out  (pivot_out_1_24),
       .r          (r_1_24)
     );

  // row 1, col 25

     reg start_in_1_25;
     wire start_out_1_25;

     reg swap_in_1_25;
     wire swap_out_1_25;

     reg [1:0] op_in_1_25;
     wire [1:0] op_out_1_25;

     wire r_1_25;

     reg data_in_1_25;
     wire data_out_1_25;

     reg pivot_in_1_25;
     wire pivot_out_1_25;

     always @(posedge clk) begin
         op_in_1_25 <= op_out_1_24;
         pivot_in_1_25 <= pivot_out_1_24;
         start_in_1_25 <= start_out_1_24;
         swap_in_1_25 <= swap_out_1_24;
     end

     always @(posedge clk) begin
         data_in_1_25 <= data_out_0_25;
     end
  
     processor_AB AB_1_25 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_25),
       .start_in   (start_in_1_25),
       .swap_in   (swap_in_1_25),
       .op_in      (op_in_1_25),
       .pivot_in   (pivot_in_1_25),
       .start_out  (start_out_1_25),
       .swap_out   (swap_out_1_25),
       .data_out   (data_out_1_25),
       .op_out     (op_out_1_25),
       .pivot_out  (pivot_out_1_25),
       .r          (r_1_25)
     );

  // row 1, col 26

     reg start_in_1_26;
     wire start_out_1_26;

     reg swap_in_1_26;
     wire swap_out_1_26;

     reg [1:0] op_in_1_26;
     wire [1:0] op_out_1_26;

     wire r_1_26;

     reg data_in_1_26;
     wire data_out_1_26;

     reg pivot_in_1_26;
     wire pivot_out_1_26;

     always @(posedge clk) begin
         op_in_1_26 <= op_out_1_25;
         pivot_in_1_26 <= pivot_out_1_25;
         start_in_1_26 <= start_out_1_25;
         swap_in_1_26 <= swap_out_1_25;
     end

     always @(posedge clk) begin
         data_in_1_26 <= data_out_0_26;
     end
  
     processor_AB AB_1_26 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_26),
       .start_in   (start_in_1_26),
       .swap_in   (swap_in_1_26),
       .op_in      (op_in_1_26),
       .pivot_in   (pivot_in_1_26),
       .start_out  (start_out_1_26),
       .swap_out   (swap_out_1_26),
       .data_out   (data_out_1_26),
       .op_out     (op_out_1_26),
       .pivot_out  (pivot_out_1_26),
       .r          (r_1_26)
     );

  // row 1, col 27

     reg start_in_1_27;
     wire start_out_1_27;

     reg swap_in_1_27;
     wire swap_out_1_27;

     reg [1:0] op_in_1_27;
     wire [1:0] op_out_1_27;

     wire r_1_27;

     reg data_in_1_27;
     wire data_out_1_27;

     reg pivot_in_1_27;
     wire pivot_out_1_27;

     always @(posedge clk) begin
         op_in_1_27 <= op_out_1_26;
         pivot_in_1_27 <= pivot_out_1_26;
         start_in_1_27 <= start_out_1_26;
         swap_in_1_27 <= swap_out_1_26;
     end

     always @(posedge clk) begin
         data_in_1_27 <= data_out_0_27;
     end
  
     processor_AB AB_1_27 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_27),
       .start_in   (start_in_1_27),
       .swap_in   (swap_in_1_27),
       .op_in      (op_in_1_27),
       .pivot_in   (pivot_in_1_27),
       .start_out  (start_out_1_27),
       .swap_out   (swap_out_1_27),
       .data_out   (data_out_1_27),
       .op_out     (op_out_1_27),
       .pivot_out  (pivot_out_1_27),
       .r          (r_1_27)
     );

  // row 1, col 28

     reg start_in_1_28;
     wire start_out_1_28;

     reg swap_in_1_28;
     wire swap_out_1_28;

     reg [1:0] op_in_1_28;
     wire [1:0] op_out_1_28;

     wire r_1_28;

     reg data_in_1_28;
     wire data_out_1_28;

     reg pivot_in_1_28;
     wire pivot_out_1_28;

     always @(posedge clk) begin
         op_in_1_28 <= op_out_1_27;
         pivot_in_1_28 <= pivot_out_1_27;
         start_in_1_28 <= start_out_1_27;
         swap_in_1_28 <= swap_out_1_27;
     end

     always @(posedge clk) begin
         data_in_1_28 <= data_out_0_28;
     end
  
     processor_AB AB_1_28 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_28),
       .start_in   (start_in_1_28),
       .swap_in   (swap_in_1_28),
       .op_in      (op_in_1_28),
       .pivot_in   (pivot_in_1_28),
       .start_out  (start_out_1_28),
       .swap_out   (swap_out_1_28),
       .data_out   (data_out_1_28),
       .op_out     (op_out_1_28),
       .pivot_out  (pivot_out_1_28),
       .r          (r_1_28)
     );

  // row 1, col 29

     reg start_in_1_29;
     wire start_out_1_29;

     reg swap_in_1_29;
     wire swap_out_1_29;

     reg [1:0] op_in_1_29;
     wire [1:0] op_out_1_29;

     wire r_1_29;

     reg data_in_1_29;
     wire data_out_1_29;

     reg pivot_in_1_29;
     wire pivot_out_1_29;

     always @(posedge clk) begin
         op_in_1_29 <= op_out_1_28;
         pivot_in_1_29 <= pivot_out_1_28;
         start_in_1_29 <= start_out_1_28;
         swap_in_1_29 <= swap_out_1_28;
     end

     always @(posedge clk) begin
         data_in_1_29 <= data_out_0_29;
     end
  
     processor_AB AB_1_29 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_29),
       .start_in   (start_in_1_29),
       .swap_in   (swap_in_1_29),
       .op_in      (op_in_1_29),
       .pivot_in   (pivot_in_1_29),
       .start_out  (start_out_1_29),
       .swap_out   (swap_out_1_29),
       .data_out   (data_out_1_29),
       .op_out     (op_out_1_29),
       .pivot_out  (pivot_out_1_29),
       .r          (r_1_29)
     );

  // row 1, col 30

     reg start_in_1_30;
     wire start_out_1_30;

     reg swap_in_1_30;
     wire swap_out_1_30;

     reg [1:0] op_in_1_30;
     wire [1:0] op_out_1_30;

     wire r_1_30;

     reg data_in_1_30;
     wire data_out_1_30;

     reg pivot_in_1_30;
     wire pivot_out_1_30;

     always @(posedge clk) begin
         op_in_1_30 <= op_out_1_29;
         pivot_in_1_30 <= pivot_out_1_29;
         start_in_1_30 <= start_out_1_29;
         swap_in_1_30 <= swap_out_1_29;
     end

     always @(posedge clk) begin
         data_in_1_30 <= data_out_0_30;
     end
  
     processor_AB AB_1_30 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_30),
       .start_in   (start_in_1_30),
       .swap_in   (swap_in_1_30),
       .op_in      (op_in_1_30),
       .pivot_in   (pivot_in_1_30),
       .start_out  (start_out_1_30),
       .swap_out   (swap_out_1_30),
       .data_out   (data_out_1_30),
       .op_out     (op_out_1_30),
       .pivot_out  (pivot_out_1_30),
       .r          (r_1_30)
     );

  // row 1, col 31

     reg start_in_1_31;
     wire start_out_1_31;

     reg swap_in_1_31;
     wire swap_out_1_31;

     reg [1:0] op_in_1_31;
     wire [1:0] op_out_1_31;

     wire r_1_31;

     reg data_in_1_31;
     wire data_out_1_31;

     reg pivot_in_1_31;
     wire pivot_out_1_31;

     always @(posedge clk) begin
         op_in_1_31 <= op_out_1_30;
         pivot_in_1_31 <= pivot_out_1_30;
         start_in_1_31 <= start_out_1_30;
         swap_in_1_31 <= swap_out_1_30;
     end

     always @(posedge clk) begin
         data_in_1_31 <= data_out_0_31;
     end
  
     processor_AB AB_1_31 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_31),
       .start_in   (start_in_1_31),
       .swap_in   (swap_in_1_31),
       .op_in      (op_in_1_31),
       .pivot_in   (pivot_in_1_31),
       .start_out  (start_out_1_31),
       .swap_out   (swap_out_1_31),
       .data_out   (data_out_1_31),
       .op_out     (op_out_1_31),
       .pivot_out  (pivot_out_1_31),
       .r          (r_1_31)
     );

  // row 1, col 32

     reg start_in_1_32;
     wire start_out_1_32;

     reg swap_in_1_32;
     wire swap_out_1_32;

     reg [1:0] op_in_1_32;
     wire [1:0] op_out_1_32;

     wire r_1_32;

     reg data_in_1_32;
     wire data_out_1_32;

     reg pivot_in_1_32;
     wire pivot_out_1_32;

     always @(posedge clk) begin
         op_in_1_32 <= op_out_1_31;
         pivot_in_1_32 <= pivot_out_1_31;
         start_in_1_32 <= start_out_1_31;
         swap_in_1_32 <= swap_out_1_31;
     end

     always @(posedge clk) begin
         data_in_1_32 <= data_out_0_32;
     end
  
     processor_AB AB_1_32 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_32),
       .start_in   (start_in_1_32),
       .swap_in   (swap_in_1_32),
       .op_in      (op_in_1_32),
       .pivot_in   (pivot_in_1_32),
       .start_out  (start_out_1_32),
       .swap_out   (swap_out_1_32),
       .data_out   (data_out_1_32),
       .op_out     (op_out_1_32),
       .pivot_out  (pivot_out_1_32),
       .r          (r_1_32)
     );

  // row 1, col 33

     reg start_in_1_33;
     wire start_out_1_33;

     reg swap_in_1_33;
     wire swap_out_1_33;

     reg [1:0] op_in_1_33;
     wire [1:0] op_out_1_33;

     wire r_1_33;

     reg data_in_1_33;
     wire data_out_1_33;

     reg pivot_in_1_33;
     wire pivot_out_1_33;

     always @(posedge clk) begin
         op_in_1_33 <= op_out_1_32;
         pivot_in_1_33 <= pivot_out_1_32;
         start_in_1_33 <= start_out_1_32;
         swap_in_1_33 <= swap_out_1_32;
     end

     always @(posedge clk) begin
         data_in_1_33 <= data_out_0_33;
     end
  
     processor_AB AB_1_33 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_33),
       .start_in   (start_in_1_33),
       .swap_in   (swap_in_1_33),
       .op_in      (op_in_1_33),
       .pivot_in   (pivot_in_1_33),
       .start_out  (start_out_1_33),
       .swap_out   (swap_out_1_33),
       .data_out   (data_out_1_33),
       .op_out     (op_out_1_33),
       .pivot_out  (pivot_out_1_33),
       .r          (r_1_33)
     );

  // row 1, col 34

     reg start_in_1_34;
     wire start_out_1_34;

     reg swap_in_1_34;
     wire swap_out_1_34;

     reg [1:0] op_in_1_34;
     wire [1:0] op_out_1_34;

     wire r_1_34;

     reg data_in_1_34;
     wire data_out_1_34;

     reg pivot_in_1_34;
     wire pivot_out_1_34;

     always @(posedge clk) begin
         op_in_1_34 <= op_out_1_33;
         pivot_in_1_34 <= pivot_out_1_33;
         start_in_1_34 <= start_out_1_33;
         swap_in_1_34 <= swap_out_1_33;
     end

     always @(posedge clk) begin
         data_in_1_34 <= data_out_0_34;
     end
  
     processor_AB AB_1_34 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_34),
       .start_in   (start_in_1_34),
       .swap_in   (swap_in_1_34),
       .op_in      (op_in_1_34),
       .pivot_in   (pivot_in_1_34),
       .start_out  (start_out_1_34),
       .swap_out   (swap_out_1_34),
       .data_out   (data_out_1_34),
       .op_out     (op_out_1_34),
       .pivot_out  (pivot_out_1_34),
       .r          (r_1_34)
     );

  // row 1, col 35

     reg start_in_1_35;
     wire start_out_1_35;

     reg swap_in_1_35;
     wire swap_out_1_35;

     reg [1:0] op_in_1_35;
     wire [1:0] op_out_1_35;

     wire r_1_35;

     reg data_in_1_35;
     wire data_out_1_35;

     reg pivot_in_1_35;
     wire pivot_out_1_35;

     always @(posedge clk) begin
         op_in_1_35 <= op_out_1_34;
         pivot_in_1_35 <= pivot_out_1_34;
         start_in_1_35 <= start_out_1_34;
         swap_in_1_35 <= swap_out_1_34;
     end

     always @(posedge clk) begin
         data_in_1_35 <= data_out_0_35;
     end
  
     processor_AB AB_1_35 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_35),
       .start_in   (start_in_1_35),
       .swap_in   (swap_in_1_35),
       .op_in      (op_in_1_35),
       .pivot_in   (pivot_in_1_35),
       .start_out  (start_out_1_35),
       .swap_out   (swap_out_1_35),
       .data_out   (data_out_1_35),
       .op_out     (op_out_1_35),
       .pivot_out  (pivot_out_1_35),
       .r          (r_1_35)
     );

  // row 1, col 36

     reg start_in_1_36;
     wire start_out_1_36;

     reg swap_in_1_36;
     wire swap_out_1_36;

     reg [1:0] op_in_1_36;
     wire [1:0] op_out_1_36;

     wire r_1_36;

     reg data_in_1_36;
     wire data_out_1_36;

     reg pivot_in_1_36;
     wire pivot_out_1_36;

     always @(posedge clk) begin
         op_in_1_36 <= op_out_1_35;
         pivot_in_1_36 <= pivot_out_1_35;
         start_in_1_36 <= start_out_1_35;
         swap_in_1_36 <= swap_out_1_35;
     end

     always @(posedge clk) begin
         data_in_1_36 <= data_out_0_36;
     end
  
     processor_AB AB_1_36 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_36),
       .start_in   (start_in_1_36),
       .swap_in   (swap_in_1_36),
       .op_in      (op_in_1_36),
       .pivot_in   (pivot_in_1_36),
       .start_out  (start_out_1_36),
       .swap_out   (swap_out_1_36),
       .data_out   (data_out_1_36),
       .op_out     (op_out_1_36),
       .pivot_out  (pivot_out_1_36),
       .r          (r_1_36)
     );

  // row 1, col 37

     reg start_in_1_37;
     wire start_out_1_37;

     reg swap_in_1_37;
     wire swap_out_1_37;

     reg [1:0] op_in_1_37;
     wire [1:0] op_out_1_37;

     wire r_1_37;

     reg data_in_1_37;
     wire data_out_1_37;

     reg pivot_in_1_37;
     wire pivot_out_1_37;

     always @(posedge clk) begin
         op_in_1_37 <= op_out_1_36;
         pivot_in_1_37 <= pivot_out_1_36;
         start_in_1_37 <= start_out_1_36;
         swap_in_1_37 <= swap_out_1_36;
     end

     always @(posedge clk) begin
         data_in_1_37 <= data_out_0_37;
     end
  
     processor_AB AB_1_37 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_37),
       .start_in   (start_in_1_37),
       .swap_in   (swap_in_1_37),
       .op_in      (op_in_1_37),
       .pivot_in   (pivot_in_1_37),
       .start_out  (start_out_1_37),
       .swap_out   (swap_out_1_37),
       .data_out   (data_out_1_37),
       .op_out     (op_out_1_37),
       .pivot_out  (pivot_out_1_37),
       .r          (r_1_37)
     );

  // row 1, col 38

     reg start_in_1_38;
     wire start_out_1_38;

     reg swap_in_1_38;
     wire swap_out_1_38;

     reg [1:0] op_in_1_38;
     wire [1:0] op_out_1_38;

     wire r_1_38;

     reg data_in_1_38;
     wire data_out_1_38;

     reg pivot_in_1_38;
     wire pivot_out_1_38;

     always @(posedge clk) begin
         op_in_1_38 <= op_out_1_37;
         pivot_in_1_38 <= pivot_out_1_37;
         start_in_1_38 <= start_out_1_37;
         swap_in_1_38 <= swap_out_1_37;
     end

     always @(posedge clk) begin
         data_in_1_38 <= data_out_0_38;
     end
  
     processor_AB AB_1_38 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_38),
       .start_in   (start_in_1_38),
       .swap_in   (swap_in_1_38),
       .op_in      (op_in_1_38),
       .pivot_in   (pivot_in_1_38),
       .start_out  (start_out_1_38),
       .swap_out   (swap_out_1_38),
       .data_out   (data_out_1_38),
       .op_out     (op_out_1_38),
       .pivot_out  (pivot_out_1_38),
       .r          (r_1_38)
     );

  // row 1, col 39

     reg start_in_1_39;
     wire start_out_1_39;

     reg swap_in_1_39;
     wire swap_out_1_39;

     reg [1:0] op_in_1_39;
     wire [1:0] op_out_1_39;

     wire r_1_39;

     reg data_in_1_39;
     wire data_out_1_39;

     reg pivot_in_1_39;
     wire pivot_out_1_39;

     always @(posedge clk) begin
         op_in_1_39 <= op_out_1_38;
         pivot_in_1_39 <= pivot_out_1_38;
         start_in_1_39 <= start_out_1_38;
         swap_in_1_39 <= swap_out_1_38;
     end

     always @(posedge clk) begin
         data_in_1_39 <= data_out_0_39;
     end
  
     processor_AB AB_1_39 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_39),
       .start_in   (start_in_1_39),
       .swap_in   (swap_in_1_39),
       .op_in      (op_in_1_39),
       .pivot_in   (pivot_in_1_39),
       .start_out  (start_out_1_39),
       .swap_out   (swap_out_1_39),
       .data_out   (data_out_1_39),
       .op_out     (op_out_1_39),
       .pivot_out  (pivot_out_1_39),
       .r          (r_1_39)
     );

  // row 1, col 40

     reg start_in_1_40;
     wire start_out_1_40;

     reg swap_in_1_40;
     wire swap_out_1_40;

     reg [1:0] op_in_1_40;
     wire [1:0] op_out_1_40;

     wire r_1_40;

     reg data_in_1_40;
     wire data_out_1_40;

     reg pivot_in_1_40;
     wire pivot_out_1_40;

     always @(posedge clk) begin
         op_in_1_40 <= op_out_1_39;
         pivot_in_1_40 <= pivot_out_1_39;
         start_in_1_40 <= start_out_1_39;
         swap_in_1_40 <= swap_out_1_39;
     end

     always @(posedge clk) begin
         data_in_1_40 <= data_out_0_40;
     end
  
     processor_AB AB_1_40 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_40),
       .start_in   (start_in_1_40),
       .swap_in   (swap_in_1_40),
       .op_in      (op_in_1_40),
       .pivot_in   (pivot_in_1_40),
       .start_out  (start_out_1_40),
       .swap_out   (swap_out_1_40),
       .data_out   (data_out_1_40),
       .op_out     (op_out_1_40),
       .pivot_out  (pivot_out_1_40),
       .r          (r_1_40)
     );

  // row 1, col 41

     reg start_in_1_41;
     wire start_out_1_41;

     reg swap_in_1_41;
     wire swap_out_1_41;

     reg [1:0] op_in_1_41;
     wire [1:0] op_out_1_41;

     wire r_1_41;

     reg data_in_1_41;
     wire data_out_1_41;

     reg pivot_in_1_41;
     wire pivot_out_1_41;

     always @(posedge clk) begin
         op_in_1_41 <= op_out_1_40;
         pivot_in_1_41 <= pivot_out_1_40;
         start_in_1_41 <= start_out_1_40;
         swap_in_1_41 <= swap_out_1_40;
     end

     always @(posedge clk) begin
         data_in_1_41 <= data_out_0_41;
     end
  
     processor_AB AB_1_41 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_41),
       .start_in   (start_in_1_41),
       .swap_in   (swap_in_1_41),
       .op_in      (op_in_1_41),
       .pivot_in   (pivot_in_1_41),
       .start_out  (start_out_1_41),
       .swap_out   (swap_out_1_41),
       .data_out   (data_out_1_41),
       .op_out     (op_out_1_41),
       .pivot_out  (pivot_out_1_41),
       .r          (r_1_41)
     );

  // row 1, col 42

     reg start_in_1_42;
     wire start_out_1_42;

     reg swap_in_1_42;
     wire swap_out_1_42;

     reg [1:0] op_in_1_42;
     wire [1:0] op_out_1_42;

     wire r_1_42;

     reg data_in_1_42;
     wire data_out_1_42;

     reg pivot_in_1_42;
     wire pivot_out_1_42;

     always @(posedge clk) begin
         op_in_1_42 <= op_out_1_41;
         pivot_in_1_42 <= pivot_out_1_41;
         start_in_1_42 <= start_out_1_41;
         swap_in_1_42 <= swap_out_1_41;
     end

     always @(posedge clk) begin
         data_in_1_42 <= data_out_0_42;
     end
  
     processor_AB AB_1_42 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_42),
       .start_in   (start_in_1_42),
       .swap_in   (swap_in_1_42),
       .op_in      (op_in_1_42),
       .pivot_in   (pivot_in_1_42),
       .start_out  (start_out_1_42),
       .swap_out   (swap_out_1_42),
       .data_out   (data_out_1_42),
       .op_out     (op_out_1_42),
       .pivot_out  (pivot_out_1_42),
       .r          (r_1_42)
     );

  // row 1, col 43

     reg start_in_1_43;
     wire start_out_1_43;

     reg swap_in_1_43;
     wire swap_out_1_43;

     reg [1:0] op_in_1_43;
     wire [1:0] op_out_1_43;

     wire r_1_43;

     reg data_in_1_43;
     wire data_out_1_43;

     reg pivot_in_1_43;
     wire pivot_out_1_43;

     always @(posedge clk) begin
         op_in_1_43 <= op_out_1_42;
         pivot_in_1_43 <= pivot_out_1_42;
         start_in_1_43 <= start_out_1_42;
         swap_in_1_43 <= swap_out_1_42;
     end

     always @(posedge clk) begin
         data_in_1_43 <= data_out_0_43;
     end
  
     processor_AB AB_1_43 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_43),
       .start_in   (start_in_1_43),
       .swap_in   (swap_in_1_43),
       .op_in      (op_in_1_43),
       .pivot_in   (pivot_in_1_43),
       .start_out  (start_out_1_43),
       .swap_out   (swap_out_1_43),
       .data_out   (data_out_1_43),
       .op_out     (op_out_1_43),
       .pivot_out  (pivot_out_1_43),
       .r          (r_1_43)
     );

  // row 1, col 44

     reg start_in_1_44;
     wire start_out_1_44;

     reg swap_in_1_44;
     wire swap_out_1_44;

     reg [1:0] op_in_1_44;
     wire [1:0] op_out_1_44;

     wire r_1_44;

     reg data_in_1_44;
     wire data_out_1_44;

     reg pivot_in_1_44;
     wire pivot_out_1_44;

     always @(posedge clk) begin
         op_in_1_44 <= op_out_1_43;
         pivot_in_1_44 <= pivot_out_1_43;
         start_in_1_44 <= start_out_1_43;
         swap_in_1_44 <= swap_out_1_43;
     end

     always @(posedge clk) begin
         data_in_1_44 <= data_out_0_44;
     end
  
     processor_AB AB_1_44 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_44),
       .start_in   (start_in_1_44),
       .swap_in   (swap_in_1_44),
       .op_in      (op_in_1_44),
       .pivot_in   (pivot_in_1_44),
       .start_out  (start_out_1_44),
       .swap_out   (swap_out_1_44),
       .data_out   (data_out_1_44),
       .op_out     (op_out_1_44),
       .pivot_out  (pivot_out_1_44),
       .r          (r_1_44)
     );

  // row 1, col 45

     reg start_in_1_45;
     wire start_out_1_45;

     reg swap_in_1_45;
     wire swap_out_1_45;

     reg [1:0] op_in_1_45;
     wire [1:0] op_out_1_45;

     wire r_1_45;

     reg data_in_1_45;
     wire data_out_1_45;

     reg pivot_in_1_45;
     wire pivot_out_1_45;

     always @(posedge clk) begin
         op_in_1_45 <= op_out_1_44;
         pivot_in_1_45 <= pivot_out_1_44;
         start_in_1_45 <= start_out_1_44;
         swap_in_1_45 <= swap_out_1_44;
     end

     always @(posedge clk) begin
         data_in_1_45 <= data_out_0_45;
     end
  
     processor_AB AB_1_45 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_45),
       .start_in   (start_in_1_45),
       .swap_in   (swap_in_1_45),
       .op_in      (op_in_1_45),
       .pivot_in   (pivot_in_1_45),
       .start_out  (start_out_1_45),
       .swap_out   (swap_out_1_45),
       .data_out   (data_out_1_45),
       .op_out     (op_out_1_45),
       .pivot_out  (pivot_out_1_45),
       .r          (r_1_45)
     );

  // row 1, col 46

     reg start_in_1_46;
     wire start_out_1_46;

     reg swap_in_1_46;
     wire swap_out_1_46;

     reg [1:0] op_in_1_46;
     wire [1:0] op_out_1_46;

     wire r_1_46;

     reg data_in_1_46;
     wire data_out_1_46;

     reg pivot_in_1_46;
     wire pivot_out_1_46;

     always @(posedge clk) begin
         op_in_1_46 <= op_out_1_45;
         pivot_in_1_46 <= pivot_out_1_45;
         start_in_1_46 <= start_out_1_45;
         swap_in_1_46 <= swap_out_1_45;
     end

     always @(posedge clk) begin
         data_in_1_46 <= data_out_0_46;
     end
  
     processor_AB AB_1_46 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_46),
       .start_in   (start_in_1_46),
       .swap_in   (swap_in_1_46),
       .op_in      (op_in_1_46),
       .pivot_in   (pivot_in_1_46),
       .start_out  (start_out_1_46),
       .swap_out   (swap_out_1_46),
       .data_out   (data_out_1_46),
       .op_out     (op_out_1_46),
       .pivot_out  (pivot_out_1_46),
       .r          (r_1_46)
     );

  // row 1, col 47

     reg start_in_1_47;
     wire start_out_1_47;

     reg swap_in_1_47;
     wire swap_out_1_47;

     reg [1:0] op_in_1_47;
     wire [1:0] op_out_1_47;

     wire r_1_47;

     reg data_in_1_47;
     wire data_out_1_47;

     reg pivot_in_1_47;
     wire pivot_out_1_47;

     always @(posedge clk) begin
         op_in_1_47 <= op_out_1_46;
         pivot_in_1_47 <= pivot_out_1_46;
         start_in_1_47 <= start_out_1_46;
         swap_in_1_47 <= swap_out_1_46;
     end

     always @(posedge clk) begin
         data_in_1_47 <= data_out_0_47;
     end
  
     processor_AB AB_1_47 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_47),
       .start_in   (start_in_1_47),
       .swap_in   (swap_in_1_47),
       .op_in      (op_in_1_47),
       .pivot_in   (pivot_in_1_47),
       .start_out  (start_out_1_47),
       .swap_out   (swap_out_1_47),
       .data_out   (data_out_1_47),
       .op_out     (op_out_1_47),
       .pivot_out  (pivot_out_1_47),
       .r          (r_1_47)
     );

  // row 1, col 48

     reg start_in_1_48;
     wire start_out_1_48;

     reg swap_in_1_48;
     wire swap_out_1_48;

     reg [1:0] op_in_1_48;
     wire [1:0] op_out_1_48;

     wire r_1_48;

     reg data_in_1_48;
     wire data_out_1_48;

     reg pivot_in_1_48;
     wire pivot_out_1_48;

     always @(posedge clk) begin
         op_in_1_48 <= op_out_1_47;
         pivot_in_1_48 <= pivot_out_1_47;
         start_in_1_48 <= start_out_1_47;
         swap_in_1_48 <= swap_out_1_47;
     end

     always @(posedge clk) begin
         data_in_1_48 <= data_out_0_48;
     end
  
     processor_AB AB_1_48 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_48),
       .start_in   (start_in_1_48),
       .swap_in   (swap_in_1_48),
       .op_in      (op_in_1_48),
       .pivot_in   (pivot_in_1_48),
       .start_out  (start_out_1_48),
       .swap_out   (swap_out_1_48),
       .data_out   (data_out_1_48),
       .op_out     (op_out_1_48),
       .pivot_out  (pivot_out_1_48),
       .r          (r_1_48)
     );

  // row 1, col 49

     reg start_in_1_49;
     wire start_out_1_49;

     reg swap_in_1_49;
     wire swap_out_1_49;

     reg [1:0] op_in_1_49;
     wire [1:0] op_out_1_49;

     wire r_1_49;

     reg data_in_1_49;
     wire data_out_1_49;

     reg pivot_in_1_49;
     wire pivot_out_1_49;

     always @(posedge clk) begin
         op_in_1_49 <= op_out_1_48;
         pivot_in_1_49 <= pivot_out_1_48;
         start_in_1_49 <= start_out_1_48;
         swap_in_1_49 <= swap_out_1_48;
     end

     always @(posedge clk) begin
         data_in_1_49 <= data_out_0_49;
     end
  
     processor_AB AB_1_49 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_49),
       .start_in   (start_in_1_49),
       .swap_in   (swap_in_1_49),
       .op_in      (op_in_1_49),
       .pivot_in   (pivot_in_1_49),
       .start_out  (start_out_1_49),
       .swap_out   (swap_out_1_49),
       .data_out   (data_out_1_49),
       .op_out     (op_out_1_49),
       .pivot_out  (pivot_out_1_49),
       .r          (r_1_49)
     );

  // row 1, col 50

     reg start_in_1_50;
     wire start_out_1_50;

     reg swap_in_1_50;
     wire swap_out_1_50;

     reg [1:0] op_in_1_50;
     wire [1:0] op_out_1_50;

     wire r_1_50;

     reg data_in_1_50;
     wire data_out_1_50;

     reg pivot_in_1_50;
     wire pivot_out_1_50;

     always @(posedge clk) begin
         op_in_1_50 <= op_out_1_49;
         pivot_in_1_50 <= pivot_out_1_49;
         start_in_1_50 <= start_out_1_49;
         swap_in_1_50 <= swap_out_1_49;
     end

     always @(posedge clk) begin
         data_in_1_50 <= data_out_0_50;
     end
  
     processor_AB AB_1_50 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_50),
       .start_in   (start_in_1_50),
       .swap_in   (swap_in_1_50),
       .op_in      (op_in_1_50),
       .pivot_in   (pivot_in_1_50),
       .start_out  (start_out_1_50),
       .swap_out   (swap_out_1_50),
       .data_out   (data_out_1_50),
       .op_out     (op_out_1_50),
       .pivot_out  (pivot_out_1_50),
       .r          (r_1_50)
     );

  // row 1, col 51

     reg start_in_1_51;
     wire start_out_1_51;

     reg swap_in_1_51;
     wire swap_out_1_51;

     reg [1:0] op_in_1_51;
     wire [1:0] op_out_1_51;

     wire r_1_51;

     reg data_in_1_51;
     wire data_out_1_51;

     reg pivot_in_1_51;
     wire pivot_out_1_51;

     always @(posedge clk) begin
         op_in_1_51 <= op_out_1_50;
         pivot_in_1_51 <= pivot_out_1_50;
         start_in_1_51 <= start_out_1_50;
         swap_in_1_51 <= swap_out_1_50;
     end

     always @(posedge clk) begin
         data_in_1_51 <= data_out_0_51;
     end
  
     processor_AB AB_1_51 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_51),
       .start_in   (start_in_1_51),
       .swap_in   (swap_in_1_51),
       .op_in      (op_in_1_51),
       .pivot_in   (pivot_in_1_51),
       .start_out  (start_out_1_51),
       .swap_out   (swap_out_1_51),
       .data_out   (data_out_1_51),
       .op_out     (op_out_1_51),
       .pivot_out  (pivot_out_1_51),
       .r          (r_1_51)
     );

  // row 1, col 52

     reg start_in_1_52;
     wire start_out_1_52;

     reg swap_in_1_52;
     wire swap_out_1_52;

     reg [1:0] op_in_1_52;
     wire [1:0] op_out_1_52;

     wire r_1_52;

     reg data_in_1_52;
     wire data_out_1_52;

     reg pivot_in_1_52;
     wire pivot_out_1_52;

     always @(posedge clk) begin
         op_in_1_52 <= op_out_1_51;
         pivot_in_1_52 <= pivot_out_1_51;
         start_in_1_52 <= start_out_1_51;
         swap_in_1_52 <= swap_out_1_51;
     end

     always @(posedge clk) begin
         data_in_1_52 <= data_out_0_52;
     end
  
     processor_AB AB_1_52 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_52),
       .start_in   (start_in_1_52),
       .swap_in   (swap_in_1_52),
       .op_in      (op_in_1_52),
       .pivot_in   (pivot_in_1_52),
       .start_out  (start_out_1_52),
       .swap_out   (swap_out_1_52),
       .data_out   (data_out_1_52),
       .op_out     (op_out_1_52),
       .pivot_out  (pivot_out_1_52),
       .r          (r_1_52)
     );

  // row 1, col 53

     reg start_in_1_53;
     wire start_out_1_53;

     reg swap_in_1_53;
     wire swap_out_1_53;

     reg [1:0] op_in_1_53;
     wire [1:0] op_out_1_53;

     wire r_1_53;

     reg data_in_1_53;
     wire data_out_1_53;

     reg pivot_in_1_53;
     wire pivot_out_1_53;

     always @(posedge clk) begin
         op_in_1_53 <= op_out_1_52;
         pivot_in_1_53 <= pivot_out_1_52;
         start_in_1_53 <= start_out_1_52;
         swap_in_1_53 <= swap_out_1_52;
     end

     always @(posedge clk) begin
         data_in_1_53 <= data_out_0_53;
     end
  
     processor_AB AB_1_53 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_53),
       .start_in   (start_in_1_53),
       .swap_in   (swap_in_1_53),
       .op_in      (op_in_1_53),
       .pivot_in   (pivot_in_1_53),
       .start_out  (start_out_1_53),
       .swap_out   (swap_out_1_53),
       .data_out   (data_out_1_53),
       .op_out     (op_out_1_53),
       .pivot_out  (pivot_out_1_53),
       .r          (r_1_53)
     );

  // row 1, col 54

     reg start_in_1_54;
     wire start_out_1_54;

     reg swap_in_1_54;
     wire swap_out_1_54;

     reg [1:0] op_in_1_54;
     wire [1:0] op_out_1_54;

     wire r_1_54;

     reg data_in_1_54;
     wire data_out_1_54;

     reg pivot_in_1_54;
     wire pivot_out_1_54;

     always @(posedge clk) begin
         op_in_1_54 <= op_out_1_53;
         pivot_in_1_54 <= pivot_out_1_53;
         start_in_1_54 <= start_out_1_53;
         swap_in_1_54 <= swap_out_1_53;
     end

     always @(posedge clk) begin
         data_in_1_54 <= data_out_0_54;
     end
  
     processor_AB AB_1_54 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_54),
       .start_in   (start_in_1_54),
       .swap_in   (swap_in_1_54),
       .op_in      (op_in_1_54),
       .pivot_in   (pivot_in_1_54),
       .start_out  (start_out_1_54),
       .swap_out   (swap_out_1_54),
       .data_out   (data_out_1_54),
       .op_out     (op_out_1_54),
       .pivot_out  (pivot_out_1_54),
       .r          (r_1_54)
     );

  // row 1, col 55

     reg start_in_1_55;
     wire start_out_1_55;

     reg swap_in_1_55;
     wire swap_out_1_55;

     reg [1:0] op_in_1_55;
     wire [1:0] op_out_1_55;

     wire r_1_55;

     reg data_in_1_55;
     wire data_out_1_55;

     reg pivot_in_1_55;
     wire pivot_out_1_55;

     always @(posedge clk) begin
         op_in_1_55 <= op_out_1_54;
         pivot_in_1_55 <= pivot_out_1_54;
         start_in_1_55 <= start_out_1_54;
         swap_in_1_55 <= swap_out_1_54;
     end

     always @(posedge clk) begin
         data_in_1_55 <= data_out_0_55;
     end
  
     processor_AB AB_1_55 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_55),
       .start_in   (start_in_1_55),
       .swap_in   (swap_in_1_55),
       .op_in      (op_in_1_55),
       .pivot_in   (pivot_in_1_55),
       .start_out  (start_out_1_55),
       .swap_out   (swap_out_1_55),
       .data_out   (data_out_1_55),
       .op_out     (op_out_1_55),
       .pivot_out  (pivot_out_1_55),
       .r          (r_1_55)
     );

  // row 1, col 56

     reg start_in_1_56;
     wire start_out_1_56;

     reg swap_in_1_56;
     wire swap_out_1_56;

     reg [1:0] op_in_1_56;
     wire [1:0] op_out_1_56;

     wire r_1_56;

     reg data_in_1_56;
     wire data_out_1_56;

     reg pivot_in_1_56;
     wire pivot_out_1_56;

     always @(posedge clk) begin
         op_in_1_56 <= op_out_1_55;
         pivot_in_1_56 <= pivot_out_1_55;
         start_in_1_56 <= start_out_1_55;
         swap_in_1_56 <= swap_out_1_55;
     end

     always @(posedge clk) begin
         data_in_1_56 <= data_out_0_56;
     end
  
     processor_AB AB_1_56 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_56),
       .start_in   (start_in_1_56),
       .swap_in   (swap_in_1_56),
       .op_in      (op_in_1_56),
       .pivot_in   (pivot_in_1_56),
       .start_out  (start_out_1_56),
       .swap_out   (swap_out_1_56),
       .data_out   (data_out_1_56),
       .op_out     (op_out_1_56),
       .pivot_out  (pivot_out_1_56),
       .r          (r_1_56)
     );

  // row 1, col 57

     reg start_in_1_57;
     wire start_out_1_57;

     reg swap_in_1_57;
     wire swap_out_1_57;

     reg [1:0] op_in_1_57;
     wire [1:0] op_out_1_57;

     wire r_1_57;

     reg data_in_1_57;
     wire data_out_1_57;

     reg pivot_in_1_57;
     wire pivot_out_1_57;

     always @(posedge clk) begin
         op_in_1_57 <= op_out_1_56;
         pivot_in_1_57 <= pivot_out_1_56;
         start_in_1_57 <= start_out_1_56;
         swap_in_1_57 <= swap_out_1_56;
     end

     always @(posedge clk) begin
         data_in_1_57 <= data_out_0_57;
     end
  
     processor_AB AB_1_57 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_57),
       .start_in   (start_in_1_57),
       .swap_in   (swap_in_1_57),
       .op_in      (op_in_1_57),
       .pivot_in   (pivot_in_1_57),
       .start_out  (start_out_1_57),
       .swap_out   (swap_out_1_57),
       .data_out   (data_out_1_57),
       .op_out     (op_out_1_57),
       .pivot_out  (pivot_out_1_57),
       .r          (r_1_57)
     );

  // row 1, col 58

     reg start_in_1_58;
     wire start_out_1_58;

     reg swap_in_1_58;
     wire swap_out_1_58;

     reg [1:0] op_in_1_58;
     wire [1:0] op_out_1_58;

     wire r_1_58;

     reg data_in_1_58;
     wire data_out_1_58;

     reg pivot_in_1_58;
     wire pivot_out_1_58;

     always @(posedge clk) begin
         op_in_1_58 <= op_out_1_57;
         pivot_in_1_58 <= pivot_out_1_57;
         start_in_1_58 <= start_out_1_57;
         swap_in_1_58 <= swap_out_1_57;
     end

     always @(posedge clk) begin
         data_in_1_58 <= data_out_0_58;
     end
  
     processor_AB AB_1_58 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_58),
       .start_in   (start_in_1_58),
       .swap_in   (swap_in_1_58),
       .op_in      (op_in_1_58),
       .pivot_in   (pivot_in_1_58),
       .start_out  (start_out_1_58),
       .swap_out   (swap_out_1_58),
       .data_out   (data_out_1_58),
       .op_out     (op_out_1_58),
       .pivot_out  (pivot_out_1_58),
       .r          (r_1_58)
     );

  // row 1, col 59

     reg start_in_1_59;
     wire start_out_1_59;

     reg swap_in_1_59;
     wire swap_out_1_59;

     reg [1:0] op_in_1_59;
     wire [1:0] op_out_1_59;

     wire r_1_59;

     reg data_in_1_59;
     wire data_out_1_59;

     reg pivot_in_1_59;
     wire pivot_out_1_59;

     always @(posedge clk) begin
         op_in_1_59 <= op_out_1_58;
         pivot_in_1_59 <= pivot_out_1_58;
         start_in_1_59 <= start_out_1_58;
         swap_in_1_59 <= swap_out_1_58;
     end

     always @(posedge clk) begin
         data_in_1_59 <= data_out_0_59;
     end
  
     processor_AB AB_1_59 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_59),
       .start_in   (start_in_1_59),
       .swap_in   (swap_in_1_59),
       .op_in      (op_in_1_59),
       .pivot_in   (pivot_in_1_59),
       .start_out  (start_out_1_59),
       .swap_out   (swap_out_1_59),
       .data_out   (data_out_1_59),
       .op_out     (op_out_1_59),
       .pivot_out  (pivot_out_1_59),
       .r          (r_1_59)
     );

  // row 1, col 60

     reg start_in_1_60;
     wire start_out_1_60;

     reg swap_in_1_60;
     wire swap_out_1_60;

     reg [1:0] op_in_1_60;
     wire [1:0] op_out_1_60;

     wire r_1_60;

     reg data_in_1_60;
     wire data_out_1_60;

     reg pivot_in_1_60;
     wire pivot_out_1_60;

     always @(posedge clk) begin
         op_in_1_60 <= op_out_1_59;
         pivot_in_1_60 <= pivot_out_1_59;
         start_in_1_60 <= start_out_1_59;
         swap_in_1_60 <= swap_out_1_59;
     end

     always @(posedge clk) begin
         data_in_1_60 <= data_out_0_60;
     end
  
     processor_AB AB_1_60 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_60),
       .start_in   (start_in_1_60),
       .swap_in   (swap_in_1_60),
       .op_in      (op_in_1_60),
       .pivot_in   (pivot_in_1_60),
       .start_out  (start_out_1_60),
       .swap_out   (swap_out_1_60),
       .data_out   (data_out_1_60),
       .op_out     (op_out_1_60),
       .pivot_out  (pivot_out_1_60),
       .r          (r_1_60)
     );

  // row 1, col 61

     reg start_in_1_61;
     wire start_out_1_61;

     reg swap_in_1_61;
     wire swap_out_1_61;

     reg [1:0] op_in_1_61;
     wire [1:0] op_out_1_61;

     wire r_1_61;

     reg data_in_1_61;
     wire data_out_1_61;

     reg pivot_in_1_61;
     wire pivot_out_1_61;

     always @(posedge clk) begin
         op_in_1_61 <= op_out_1_60;
         pivot_in_1_61 <= pivot_out_1_60;
         start_in_1_61 <= start_out_1_60;
         swap_in_1_61 <= swap_out_1_60;
     end

     always @(posedge clk) begin
         data_in_1_61 <= data_out_0_61;
     end
  
     processor_AB AB_1_61 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_61),
       .start_in   (start_in_1_61),
       .swap_in   (swap_in_1_61),
       .op_in      (op_in_1_61),
       .pivot_in   (pivot_in_1_61),
       .start_out  (start_out_1_61),
       .swap_out   (swap_out_1_61),
       .data_out   (data_out_1_61),
       .op_out     (op_out_1_61),
       .pivot_out  (pivot_out_1_61),
       .r          (r_1_61)
     );

  // row 1, col 62

     reg start_in_1_62;
     wire start_out_1_62;

     reg swap_in_1_62;
     wire swap_out_1_62;

     reg [1:0] op_in_1_62;
     wire [1:0] op_out_1_62;

     wire r_1_62;

     reg data_in_1_62;
     wire data_out_1_62;

     reg pivot_in_1_62;
     wire pivot_out_1_62;

     always @(posedge clk) begin
         op_in_1_62 <= op_out_1_61;
         pivot_in_1_62 <= pivot_out_1_61;
         start_in_1_62 <= start_out_1_61;
         swap_in_1_62 <= swap_out_1_61;
     end

     always @(posedge clk) begin
         data_in_1_62 <= data_out_0_62;
     end
  
     processor_AB AB_1_62 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_62),
       .start_in   (start_in_1_62),
       .swap_in   (swap_in_1_62),
       .op_in      (op_in_1_62),
       .pivot_in   (pivot_in_1_62),
       .start_out  (start_out_1_62),
       .swap_out   (swap_out_1_62),
       .data_out   (data_out_1_62),
       .op_out     (op_out_1_62),
       .pivot_out  (pivot_out_1_62),
       .r          (r_1_62)
     );

  // row 1, col 63

     reg start_in_1_63;
     wire start_out_1_63;

     reg swap_in_1_63;
     wire swap_out_1_63;

     reg [1:0] op_in_1_63;
     wire [1:0] op_out_1_63;

     wire r_1_63;

     reg data_in_1_63;
     wire data_out_1_63;

     reg pivot_in_1_63;
     wire pivot_out_1_63;

     always @(posedge clk) begin
         op_in_1_63 <= op_out_1_62;
         pivot_in_1_63 <= pivot_out_1_62;
         start_in_1_63 <= start_out_1_62;
         swap_in_1_63 <= swap_out_1_62;
     end

     always @(posedge clk) begin
         data_in_1_63 <= data_out_0_63;
     end
  
     processor_AB AB_1_63 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_63),
       .start_in   (start_in_1_63),
       .swap_in   (swap_in_1_63),
       .op_in      (op_in_1_63),
       .pivot_in   (pivot_in_1_63),
       .start_out  (start_out_1_63),
       .swap_out   (swap_out_1_63),
       .data_out   (data_out_1_63),
       .op_out     (op_out_1_63),
       .pivot_out  (pivot_out_1_63),
       .r          (r_1_63)
     );

  // row 1, col 64

     reg start_in_1_64;
     wire start_out_1_64;

     reg swap_in_1_64;
     wire swap_out_1_64;

     reg [1:0] op_in_1_64;
     wire [1:0] op_out_1_64;

     wire r_1_64;

     reg data_in_1_64;
     wire data_out_1_64;

     reg pivot_in_1_64;
     wire pivot_out_1_64;

     always @(posedge clk) begin
         op_in_1_64 <= op_out_1_63;
         pivot_in_1_64 <= pivot_out_1_63;
         start_in_1_64 <= start_out_1_63;
         swap_in_1_64 <= swap_out_1_63;
     end

     always @(posedge clk) begin
         data_in_1_64 <= data_out_0_64;
     end
  
     processor_AB AB_1_64 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_64),
       .start_in   (start_in_1_64),
       .swap_in   (swap_in_1_64),
       .op_in      (op_in_1_64),
       .pivot_in   (pivot_in_1_64),
       .start_out  (start_out_1_64),
       .swap_out   (swap_out_1_64),
       .data_out   (data_out_1_64),
       .op_out     (op_out_1_64),
       .pivot_out  (pivot_out_1_64),
       .r          (r_1_64)
     );

  // row 1, col 65

     reg start_in_1_65;
     wire start_out_1_65;

     reg swap_in_1_65;
     wire swap_out_1_65;

     reg [1:0] op_in_1_65;
     wire [1:0] op_out_1_65;

     wire r_1_65;

     reg data_in_1_65;
     wire data_out_1_65;

     reg pivot_in_1_65;
     wire pivot_out_1_65;

     always @(posedge clk) begin
         op_in_1_65 <= op_out_1_64;
         pivot_in_1_65 <= pivot_out_1_64;
         start_in_1_65 <= start_out_1_64;
         swap_in_1_65 <= swap_out_1_64;
     end

     always @(posedge clk) begin
         data_in_1_65 <= data_out_0_65;
     end
  
     processor_AB AB_1_65 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_65),
       .start_in   (start_in_1_65),
       .swap_in   (swap_in_1_65),
       .op_in      (op_in_1_65),
       .pivot_in   (pivot_in_1_65),
       .start_out  (start_out_1_65),
       .swap_out   (swap_out_1_65),
       .data_out   (data_out_1_65),
       .op_out     (op_out_1_65),
       .pivot_out  (pivot_out_1_65),
       .r          (r_1_65)
     );

  // row 1, col 66

     reg start_in_1_66;
     wire start_out_1_66;

     reg swap_in_1_66;
     wire swap_out_1_66;

     reg [1:0] op_in_1_66;
     wire [1:0] op_out_1_66;

     wire r_1_66;

     reg data_in_1_66;
     wire data_out_1_66;

     reg pivot_in_1_66;
     wire pivot_out_1_66;

     always @(posedge clk) begin
         op_in_1_66 <= op_out_1_65;
         pivot_in_1_66 <= pivot_out_1_65;
         start_in_1_66 <= start_out_1_65;
         swap_in_1_66 <= swap_out_1_65;
     end

     always @(posedge clk) begin
         data_in_1_66 <= data_out_0_66;
     end
  
     processor_AB AB_1_66 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_66),
       .start_in   (start_in_1_66),
       .swap_in   (swap_in_1_66),
       .op_in      (op_in_1_66),
       .pivot_in   (pivot_in_1_66),
       .start_out  (start_out_1_66),
       .swap_out   (swap_out_1_66),
       .data_out   (data_out_1_66),
       .op_out     (op_out_1_66),
       .pivot_out  (pivot_out_1_66),
       .r          (r_1_66)
     );

  // row 1, col 67

     reg start_in_1_67;
     wire start_out_1_67;

     reg swap_in_1_67;
     wire swap_out_1_67;

     reg [1:0] op_in_1_67;
     wire [1:0] op_out_1_67;

     wire r_1_67;

     reg data_in_1_67;
     wire data_out_1_67;

     reg pivot_in_1_67;
     wire pivot_out_1_67;

     always @(posedge clk) begin
         op_in_1_67 <= op_out_1_66;
         pivot_in_1_67 <= pivot_out_1_66;
         start_in_1_67 <= start_out_1_66;
         swap_in_1_67 <= swap_out_1_66;
     end

     always @(posedge clk) begin
         data_in_1_67 <= data_out_0_67;
     end
  
     processor_AB AB_1_67 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_67),
       .start_in   (start_in_1_67),
       .swap_in   (swap_in_1_67),
       .op_in      (op_in_1_67),
       .pivot_in   (pivot_in_1_67),
       .start_out  (start_out_1_67),
       .swap_out   (swap_out_1_67),
       .data_out   (data_out_1_67),
       .op_out     (op_out_1_67),
       .pivot_out  (pivot_out_1_67),
       .r          (r_1_67)
     );

  // row 1, col 68

     reg start_in_1_68;
     wire start_out_1_68;

     reg swap_in_1_68;
     wire swap_out_1_68;

     reg [1:0] op_in_1_68;
     wire [1:0] op_out_1_68;

     wire r_1_68;

     reg data_in_1_68;
     wire data_out_1_68;

     reg pivot_in_1_68;
     wire pivot_out_1_68;

     always @(posedge clk) begin
         op_in_1_68 <= op_out_1_67;
         pivot_in_1_68 <= pivot_out_1_67;
         start_in_1_68 <= start_out_1_67;
         swap_in_1_68 <= swap_out_1_67;
     end

     always @(posedge clk) begin
         data_in_1_68 <= data_out_0_68;
     end
  
     processor_AB AB_1_68 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_68),
       .start_in   (start_in_1_68),
       .swap_in   (swap_in_1_68),
       .op_in      (op_in_1_68),
       .pivot_in   (pivot_in_1_68),
       .start_out  (start_out_1_68),
       .swap_out   (swap_out_1_68),
       .data_out   (data_out_1_68),
       .op_out     (op_out_1_68),
       .pivot_out  (pivot_out_1_68),
       .r          (r_1_68)
     );

  // row 1, col 69

     reg start_in_1_69;
     wire start_out_1_69;

     reg swap_in_1_69;
     wire swap_out_1_69;

     reg [1:0] op_in_1_69;
     wire [1:0] op_out_1_69;

     wire r_1_69;

     reg data_in_1_69;
     wire data_out_1_69;

     reg pivot_in_1_69;
     wire pivot_out_1_69;

     always @(posedge clk) begin
         op_in_1_69 <= op_out_1_68;
         pivot_in_1_69 <= pivot_out_1_68;
         start_in_1_69 <= start_out_1_68;
         swap_in_1_69 <= swap_out_1_68;
     end

     always @(posedge clk) begin
         data_in_1_69 <= data_out_0_69;
     end
  
     processor_AB AB_1_69 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_69),
       .start_in   (start_in_1_69),
       .swap_in   (swap_in_1_69),
       .op_in      (op_in_1_69),
       .pivot_in   (pivot_in_1_69),
       .start_out  (start_out_1_69),
       .swap_out   (swap_out_1_69),
       .data_out   (data_out_1_69),
       .op_out     (op_out_1_69),
       .pivot_out  (pivot_out_1_69),
       .r          (r_1_69)
     );

  // row 1, col 70

     reg start_in_1_70;
     wire start_out_1_70;

     reg swap_in_1_70;
     wire swap_out_1_70;

     reg [1:0] op_in_1_70;
     wire [1:0] op_out_1_70;

     wire r_1_70;

     reg data_in_1_70;
     wire data_out_1_70;

     reg pivot_in_1_70;
     wire pivot_out_1_70;

     always @(posedge clk) begin
         op_in_1_70 <= op_out_1_69;
         pivot_in_1_70 <= pivot_out_1_69;
         start_in_1_70 <= start_out_1_69;
         swap_in_1_70 <= swap_out_1_69;
     end

     always @(posedge clk) begin
         data_in_1_70 <= data_out_0_70;
     end
  
     processor_AB AB_1_70 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_70),
       .start_in   (start_in_1_70),
       .swap_in   (swap_in_1_70),
       .op_in      (op_in_1_70),
       .pivot_in   (pivot_in_1_70),
       .start_out  (start_out_1_70),
       .swap_out   (swap_out_1_70),
       .data_out   (data_out_1_70),
       .op_out     (op_out_1_70),
       .pivot_out  (pivot_out_1_70),
       .r          (r_1_70)
     );

  // row 1, col 71

     reg start_in_1_71;
     wire start_out_1_71;

     reg swap_in_1_71;
     wire swap_out_1_71;

     reg [1:0] op_in_1_71;
     wire [1:0] op_out_1_71;

     wire r_1_71;

     reg data_in_1_71;
     wire data_out_1_71;

     reg pivot_in_1_71;
     wire pivot_out_1_71;

     always @(posedge clk) begin
         op_in_1_71 <= op_out_1_70;
         pivot_in_1_71 <= pivot_out_1_70;
         start_in_1_71 <= start_out_1_70;
         swap_in_1_71 <= swap_out_1_70;
     end

     always @(posedge clk) begin
         data_in_1_71 <= data_out_0_71;
     end
  
     processor_AB AB_1_71 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_71),
       .start_in   (start_in_1_71),
       .swap_in   (swap_in_1_71),
       .op_in      (op_in_1_71),
       .pivot_in   (pivot_in_1_71),
       .start_out  (start_out_1_71),
       .swap_out   (swap_out_1_71),
       .data_out   (data_out_1_71),
       .op_out     (op_out_1_71),
       .pivot_out  (pivot_out_1_71),
       .r          (r_1_71)
     );

  // row 1, col 72

     reg start_in_1_72;
     wire start_out_1_72;

     reg swap_in_1_72;
     wire swap_out_1_72;

     reg [1:0] op_in_1_72;
     wire [1:0] op_out_1_72;

     wire r_1_72;

     reg data_in_1_72;
     wire data_out_1_72;

     reg pivot_in_1_72;
     wire pivot_out_1_72;

     always @(posedge clk) begin
         op_in_1_72 <= op_out_1_71;
         pivot_in_1_72 <= pivot_out_1_71;
         start_in_1_72 <= start_out_1_71;
         swap_in_1_72 <= swap_out_1_71;
     end

     always @(posedge clk) begin
         data_in_1_72 <= data_out_0_72;
     end
  
     processor_AB AB_1_72 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_72),
       .start_in   (start_in_1_72),
       .swap_in   (swap_in_1_72),
       .op_in      (op_in_1_72),
       .pivot_in   (pivot_in_1_72),
       .start_out  (start_out_1_72),
       .swap_out   (swap_out_1_72),
       .data_out   (data_out_1_72),
       .op_out     (op_out_1_72),
       .pivot_out  (pivot_out_1_72),
       .r          (r_1_72)
     );

  // row 1, col 73

     reg start_in_1_73;
     wire start_out_1_73;

     reg swap_in_1_73;
     wire swap_out_1_73;

     reg [1:0] op_in_1_73;
     wire [1:0] op_out_1_73;

     wire r_1_73;

     reg data_in_1_73;
     wire data_out_1_73;

     reg pivot_in_1_73;
     wire pivot_out_1_73;

     always @(posedge clk) begin
         op_in_1_73 <= op_out_1_72;
         pivot_in_1_73 <= pivot_out_1_72;
         start_in_1_73 <= start_out_1_72;
         swap_in_1_73 <= swap_out_1_72;
     end

     always @(posedge clk) begin
         data_in_1_73 <= data_out_0_73;
     end
  
     processor_AB AB_1_73 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_73),
       .start_in   (start_in_1_73),
       .swap_in   (swap_in_1_73),
       .op_in      (op_in_1_73),
       .pivot_in   (pivot_in_1_73),
       .start_out  (start_out_1_73),
       .swap_out   (swap_out_1_73),
       .data_out   (data_out_1_73),
       .op_out     (op_out_1_73),
       .pivot_out  (pivot_out_1_73),
       .r          (r_1_73)
     );

  // row 1, col 74

     reg start_in_1_74;
     wire start_out_1_74;

     reg swap_in_1_74;
     wire swap_out_1_74;

     reg [1:0] op_in_1_74;
     wire [1:0] op_out_1_74;

     wire r_1_74;

     reg data_in_1_74;
     wire data_out_1_74;

     reg pivot_in_1_74;
     wire pivot_out_1_74;

     always @(posedge clk) begin
         op_in_1_74 <= op_out_1_73;
         pivot_in_1_74 <= pivot_out_1_73;
         start_in_1_74 <= start_out_1_73;
         swap_in_1_74 <= swap_out_1_73;
     end

     always @(posedge clk) begin
         data_in_1_74 <= data_out_0_74;
     end
  
     processor_AB AB_1_74 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_74),
       .start_in   (start_in_1_74),
       .swap_in   (swap_in_1_74),
       .op_in      (op_in_1_74),
       .pivot_in   (pivot_in_1_74),
       .start_out  (start_out_1_74),
       .swap_out   (swap_out_1_74),
       .data_out   (data_out_1_74),
       .op_out     (op_out_1_74),
       .pivot_out  (pivot_out_1_74),
       .r          (r_1_74)
     );

  // row 1, col 75

     reg start_in_1_75;
     wire start_out_1_75;

     reg swap_in_1_75;
     wire swap_out_1_75;

     reg [1:0] op_in_1_75;
     wire [1:0] op_out_1_75;

     wire r_1_75;

     reg data_in_1_75;
     wire data_out_1_75;

     reg pivot_in_1_75;
     wire pivot_out_1_75;

     always @(posedge clk) begin
         op_in_1_75 <= op_out_1_74;
         pivot_in_1_75 <= pivot_out_1_74;
         start_in_1_75 <= start_out_1_74;
         swap_in_1_75 <= swap_out_1_74;
     end

     always @(posedge clk) begin
         data_in_1_75 <= data_out_0_75;
     end
  
     processor_AB AB_1_75 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_75),
       .start_in   (start_in_1_75),
       .swap_in   (swap_in_1_75),
       .op_in      (op_in_1_75),
       .pivot_in   (pivot_in_1_75),
       .start_out  (start_out_1_75),
       .swap_out   (swap_out_1_75),
       .data_out   (data_out_1_75),
       .op_out     (op_out_1_75),
       .pivot_out  (pivot_out_1_75),
       .r          (r_1_75)
     );

  // row 1, col 76

     reg start_in_1_76;
     wire start_out_1_76;

     reg swap_in_1_76;
     wire swap_out_1_76;

     reg [1:0] op_in_1_76;
     wire [1:0] op_out_1_76;

     wire r_1_76;

     reg data_in_1_76;
     wire data_out_1_76;

     reg pivot_in_1_76;
     wire pivot_out_1_76;

     always @(posedge clk) begin
         op_in_1_76 <= op_out_1_75;
         pivot_in_1_76 <= pivot_out_1_75;
         start_in_1_76 <= start_out_1_75;
         swap_in_1_76 <= swap_out_1_75;
     end

     always @(posedge clk) begin
         data_in_1_76 <= data_out_0_76;
     end
  
     processor_AB AB_1_76 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_76),
       .start_in   (start_in_1_76),
       .swap_in   (swap_in_1_76),
       .op_in      (op_in_1_76),
       .pivot_in   (pivot_in_1_76),
       .start_out  (start_out_1_76),
       .swap_out   (swap_out_1_76),
       .data_out   (data_out_1_76),
       .op_out     (op_out_1_76),
       .pivot_out  (pivot_out_1_76),
       .r          (r_1_76)
     );

  // row 1, col 77

     reg start_in_1_77;
     wire start_out_1_77;

     reg swap_in_1_77;
     wire swap_out_1_77;

     reg [1:0] op_in_1_77;
     wire [1:0] op_out_1_77;

     wire r_1_77;

     reg data_in_1_77;
     wire data_out_1_77;

     reg pivot_in_1_77;
     wire pivot_out_1_77;

     always @(posedge clk) begin
         op_in_1_77 <= op_out_1_76;
         pivot_in_1_77 <= pivot_out_1_76;
         start_in_1_77 <= start_out_1_76;
         swap_in_1_77 <= swap_out_1_76;
     end

     always @(posedge clk) begin
         data_in_1_77 <= data_out_0_77;
     end
  
     processor_AB AB_1_77 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_77),
       .start_in   (start_in_1_77),
       .swap_in   (swap_in_1_77),
       .op_in      (op_in_1_77),
       .pivot_in   (pivot_in_1_77),
       .start_out  (start_out_1_77),
       .swap_out   (swap_out_1_77),
       .data_out   (data_out_1_77),
       .op_out     (op_out_1_77),
       .pivot_out  (pivot_out_1_77),
       .r          (r_1_77)
     );

  // row 1, col 78

     reg start_in_1_78;
     wire start_out_1_78;

     reg swap_in_1_78;
     wire swap_out_1_78;

     reg [1:0] op_in_1_78;
     wire [1:0] op_out_1_78;

     wire r_1_78;

     reg data_in_1_78;
     wire data_out_1_78;

     reg pivot_in_1_78;
     wire pivot_out_1_78;

     always @(posedge clk) begin
         op_in_1_78 <= op_out_1_77;
         pivot_in_1_78 <= pivot_out_1_77;
         start_in_1_78 <= start_out_1_77;
         swap_in_1_78 <= swap_out_1_77;
     end

     always @(posedge clk) begin
         data_in_1_78 <= data_out_0_78;
     end
  
     processor_AB AB_1_78 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_78),
       .start_in   (start_in_1_78),
       .swap_in   (swap_in_1_78),
       .op_in      (op_in_1_78),
       .pivot_in   (pivot_in_1_78),
       .start_out  (start_out_1_78),
       .swap_out   (swap_out_1_78),
       .data_out   (data_out_1_78),
       .op_out     (op_out_1_78),
       .pivot_out  (pivot_out_1_78),
       .r          (r_1_78)
     );

  // row 1, col 79

     reg start_in_1_79;
     wire start_out_1_79;

     reg swap_in_1_79;
     wire swap_out_1_79;

     reg [1:0] op_in_1_79;
     wire [1:0] op_out_1_79;

     wire r_1_79;

     reg data_in_1_79;
     wire data_out_1_79;

     reg pivot_in_1_79;
     wire pivot_out_1_79;

     always @(posedge clk) begin
         op_in_1_79 <= op_out_1_78;
         pivot_in_1_79 <= pivot_out_1_78;
         start_in_1_79 <= start_out_1_78;
         swap_in_1_79 <= swap_out_1_78;
     end

     always @(posedge clk) begin
         data_in_1_79 <= data_out_0_79;
     end
  
     processor_AB AB_1_79 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_79),
       .start_in   (start_in_1_79),
       .swap_in   (swap_in_1_79),
       .op_in      (op_in_1_79),
       .pivot_in   (pivot_in_1_79),
       .start_out  (start_out_1_79),
       .swap_out   (swap_out_1_79),
       .data_out   (data_out_1_79),
       .op_out     (op_out_1_79),
       .pivot_out  (pivot_out_1_79),
       .r          (r_1_79)
     );

  // row 1, col 80

     reg start_in_1_80;
     wire start_out_1_80;

     reg swap_in_1_80;
     wire swap_out_1_80;

     reg [1:0] op_in_1_80;
     wire [1:0] op_out_1_80;

     wire r_1_80;

     reg data_in_1_80;
     wire data_out_1_80;

     reg pivot_in_1_80;
     wire pivot_out_1_80;

     always @(posedge clk) begin
         op_in_1_80 <= op_out_1_79;
         pivot_in_1_80 <= pivot_out_1_79;
         start_in_1_80 <= start_out_1_79;
         swap_in_1_80 <= swap_out_1_79;
     end

     always @(posedge clk) begin
         data_in_1_80 <= data_out_0_80;
     end
  
     processor_AB AB_1_80 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_80),
       .start_in   (start_in_1_80),
       .swap_in   (swap_in_1_80),
       .op_in      (op_in_1_80),
       .pivot_in   (pivot_in_1_80),
       .start_out  (start_out_1_80),
       .swap_out   (swap_out_1_80),
       .data_out   (data_out_1_80),
       .op_out     (op_out_1_80),
       .pivot_out  (pivot_out_1_80),
       .r          (r_1_80)
     );

  // row 1, col 81

     reg start_in_1_81;
     wire start_out_1_81;

     reg swap_in_1_81;
     wire swap_out_1_81;

     reg [1:0] op_in_1_81;
     wire [1:0] op_out_1_81;

     wire r_1_81;

     reg data_in_1_81;
     wire data_out_1_81;

     reg pivot_in_1_81;
     wire pivot_out_1_81;

     always @(posedge clk) begin
         op_in_1_81 <= op_out_1_80;
         pivot_in_1_81 <= pivot_out_1_80;
         start_in_1_81 <= start_out_1_80;
         swap_in_1_81 <= swap_out_1_80;
     end

     always @(posedge clk) begin
         data_in_1_81 <= data_out_0_81;
     end
  
     processor_AB AB_1_81 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_81),
       .start_in   (start_in_1_81),
       .swap_in   (swap_in_1_81),
       .op_in      (op_in_1_81),
       .pivot_in   (pivot_in_1_81),
       .start_out  (start_out_1_81),
       .swap_out   (swap_out_1_81),
       .data_out   (data_out_1_81),
       .op_out     (op_out_1_81),
       .pivot_out  (pivot_out_1_81),
       .r          (r_1_81)
     );

  // row 1, col 82

     reg start_in_1_82;
     wire start_out_1_82;

     reg swap_in_1_82;
     wire swap_out_1_82;

     reg [1:0] op_in_1_82;
     wire [1:0] op_out_1_82;

     wire r_1_82;

     reg data_in_1_82;
     wire data_out_1_82;

     reg pivot_in_1_82;
     wire pivot_out_1_82;

     always @(posedge clk) begin
         op_in_1_82 <= op_out_1_81;
         pivot_in_1_82 <= pivot_out_1_81;
         start_in_1_82 <= start_out_1_81;
         swap_in_1_82 <= swap_out_1_81;
     end

     always @(posedge clk) begin
         data_in_1_82 <= data_out_0_82;
     end
  
     processor_AB AB_1_82 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_82),
       .start_in   (start_in_1_82),
       .swap_in   (swap_in_1_82),
       .op_in      (op_in_1_82),
       .pivot_in   (pivot_in_1_82),
       .start_out  (start_out_1_82),
       .swap_out   (swap_out_1_82),
       .data_out   (data_out_1_82),
       .op_out     (op_out_1_82),
       .pivot_out  (pivot_out_1_82),
       .r          (r_1_82)
     );

  // row 1, col 83

     reg start_in_1_83;
     wire start_out_1_83;

     reg swap_in_1_83;
     wire swap_out_1_83;

     reg [1:0] op_in_1_83;
     wire [1:0] op_out_1_83;

     wire r_1_83;

     reg data_in_1_83;
     wire data_out_1_83;

     reg pivot_in_1_83;
     wire pivot_out_1_83;

     always @(posedge clk) begin
         op_in_1_83 <= op_out_1_82;
         pivot_in_1_83 <= pivot_out_1_82;
         start_in_1_83 <= start_out_1_82;
         swap_in_1_83 <= swap_out_1_82;
     end

     always @(posedge clk) begin
         data_in_1_83 <= data_out_0_83;
     end
  
     processor_AB AB_1_83 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_83),
       .start_in   (start_in_1_83),
       .swap_in   (swap_in_1_83),
       .op_in      (op_in_1_83),
       .pivot_in   (pivot_in_1_83),
       .start_out  (start_out_1_83),
       .swap_out   (swap_out_1_83),
       .data_out   (data_out_1_83),
       .op_out     (op_out_1_83),
       .pivot_out  (pivot_out_1_83),
       .r          (r_1_83)
     );

  // row 1, col 84

     reg start_in_1_84;
     wire start_out_1_84;

     reg swap_in_1_84;
     wire swap_out_1_84;

     reg [1:0] op_in_1_84;
     wire [1:0] op_out_1_84;

     wire r_1_84;

     reg data_in_1_84;
     wire data_out_1_84;

     reg pivot_in_1_84;
     wire pivot_out_1_84;

     always @(posedge clk) begin
         op_in_1_84 <= op_out_1_83;
         pivot_in_1_84 <= pivot_out_1_83;
         start_in_1_84 <= start_out_1_83;
         swap_in_1_84 <= swap_out_1_83;
     end

     always @(posedge clk) begin
         data_in_1_84 <= data_out_0_84;
     end
  
     processor_AB AB_1_84 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_84),
       .start_in   (start_in_1_84),
       .swap_in   (swap_in_1_84),
       .op_in      (op_in_1_84),
       .pivot_in   (pivot_in_1_84),
       .start_out  (start_out_1_84),
       .swap_out   (swap_out_1_84),
       .data_out   (data_out_1_84),
       .op_out     (op_out_1_84),
       .pivot_out  (pivot_out_1_84),
       .r          (r_1_84)
     );

  // row 1, col 85

     reg start_in_1_85;
     wire start_out_1_85;

     reg swap_in_1_85;
     wire swap_out_1_85;

     reg [1:0] op_in_1_85;
     wire [1:0] op_out_1_85;

     wire r_1_85;

     reg data_in_1_85;
     wire data_out_1_85;

     reg pivot_in_1_85;
     wire pivot_out_1_85;

     always @(posedge clk) begin
         op_in_1_85 <= op_out_1_84;
         pivot_in_1_85 <= pivot_out_1_84;
         start_in_1_85 <= start_out_1_84;
         swap_in_1_85 <= swap_out_1_84;
     end

     always @(posedge clk) begin
         data_in_1_85 <= data_out_0_85;
     end
  
     processor_AB AB_1_85 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_85),
       .start_in   (start_in_1_85),
       .swap_in   (swap_in_1_85),
       .op_in      (op_in_1_85),
       .pivot_in   (pivot_in_1_85),
       .start_out  (start_out_1_85),
       .swap_out   (swap_out_1_85),
       .data_out   (data_out_1_85),
       .op_out     (op_out_1_85),
       .pivot_out  (pivot_out_1_85),
       .r          (r_1_85)
     );

  // row 1, col 86

     reg start_in_1_86;
     wire start_out_1_86;

     reg swap_in_1_86;
     wire swap_out_1_86;

     reg [1:0] op_in_1_86;
     wire [1:0] op_out_1_86;

     wire r_1_86;

     reg data_in_1_86;
     wire data_out_1_86;

     reg pivot_in_1_86;
     wire pivot_out_1_86;

     always @(posedge clk) begin
         op_in_1_86 <= op_out_1_85;
         pivot_in_1_86 <= pivot_out_1_85;
         start_in_1_86 <= start_out_1_85;
         swap_in_1_86 <= swap_out_1_85;
     end

     always @(posedge clk) begin
         data_in_1_86 <= data_out_0_86;
     end
  
     processor_AB AB_1_86 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_86),
       .start_in   (start_in_1_86),
       .swap_in   (swap_in_1_86),
       .op_in      (op_in_1_86),
       .pivot_in   (pivot_in_1_86),
       .start_out  (start_out_1_86),
       .swap_out   (swap_out_1_86),
       .data_out   (data_out_1_86),
       .op_out     (op_out_1_86),
       .pivot_out  (pivot_out_1_86),
       .r          (r_1_86)
     );

  // row 1, col 87

     reg start_in_1_87;
     wire start_out_1_87;

     reg swap_in_1_87;
     wire swap_out_1_87;

     reg [1:0] op_in_1_87;
     wire [1:0] op_out_1_87;

     wire r_1_87;

     reg data_in_1_87;
     wire data_out_1_87;

     reg pivot_in_1_87;
     wire pivot_out_1_87;

     always @(posedge clk) begin
         op_in_1_87 <= op_out_1_86;
         pivot_in_1_87 <= pivot_out_1_86;
         start_in_1_87 <= start_out_1_86;
         swap_in_1_87 <= swap_out_1_86;
     end

     always @(posedge clk) begin
         data_in_1_87 <= data_out_0_87;
     end
  
     processor_AB AB_1_87 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_87),
       .start_in   (start_in_1_87),
       .swap_in   (swap_in_1_87),
       .op_in      (op_in_1_87),
       .pivot_in   (pivot_in_1_87),
       .start_out  (start_out_1_87),
       .swap_out   (swap_out_1_87),
       .data_out   (data_out_1_87),
       .op_out     (op_out_1_87),
       .pivot_out  (pivot_out_1_87),
       .r          (r_1_87)
     );

  // row 1, col 88

     reg start_in_1_88;
     wire start_out_1_88;

     reg swap_in_1_88;
     wire swap_out_1_88;

     reg [1:0] op_in_1_88;
     wire [1:0] op_out_1_88;

     wire r_1_88;

     reg data_in_1_88;
     wire data_out_1_88;

     reg pivot_in_1_88;
     wire pivot_out_1_88;

     always @(posedge clk) begin
         op_in_1_88 <= op_out_1_87;
         pivot_in_1_88 <= pivot_out_1_87;
         start_in_1_88 <= start_out_1_87;
         swap_in_1_88 <= swap_out_1_87;
     end

     always @(posedge clk) begin
         data_in_1_88 <= data_out_0_88;
     end
  
     processor_AB AB_1_88 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_88),
       .start_in   (start_in_1_88),
       .swap_in   (swap_in_1_88),
       .op_in      (op_in_1_88),
       .pivot_in   (pivot_in_1_88),
       .start_out  (start_out_1_88),
       .swap_out   (swap_out_1_88),
       .data_out   (data_out_1_88),
       .op_out     (op_out_1_88),
       .pivot_out  (pivot_out_1_88),
       .r          (r_1_88)
     );

  // row 1, col 89

     reg start_in_1_89;
     wire start_out_1_89;

     reg swap_in_1_89;
     wire swap_out_1_89;

     reg [1:0] op_in_1_89;
     wire [1:0] op_out_1_89;

     wire r_1_89;

     reg data_in_1_89;
     wire data_out_1_89;

     reg pivot_in_1_89;
     wire pivot_out_1_89;

     always @(posedge clk) begin
         op_in_1_89 <= op_out_1_88;
         pivot_in_1_89 <= pivot_out_1_88;
         start_in_1_89 <= start_out_1_88;
         swap_in_1_89 <= swap_out_1_88;
     end

     always @(posedge clk) begin
         data_in_1_89 <= data_out_0_89;
     end
  
     processor_AB AB_1_89 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_89),
       .start_in   (start_in_1_89),
       .swap_in   (swap_in_1_89),
       .op_in      (op_in_1_89),
       .pivot_in   (pivot_in_1_89),
       .start_out  (start_out_1_89),
       .swap_out   (swap_out_1_89),
       .data_out   (data_out_1_89),
       .op_out     (op_out_1_89),
       .pivot_out  (pivot_out_1_89),
       .r          (r_1_89)
     );

  // row 1, col 90

     reg start_in_1_90;
     wire start_out_1_90;

     reg swap_in_1_90;
     wire swap_out_1_90;

     reg [1:0] op_in_1_90;
     wire [1:0] op_out_1_90;

     wire r_1_90;

     reg data_in_1_90;
     wire data_out_1_90;

     reg pivot_in_1_90;
     wire pivot_out_1_90;

     always @(posedge clk) begin
         op_in_1_90 <= op_out_1_89;
         pivot_in_1_90 <= pivot_out_1_89;
         start_in_1_90 <= start_out_1_89;
         swap_in_1_90 <= swap_out_1_89;
     end

     always @(posedge clk) begin
         data_in_1_90 <= data_out_0_90;
     end
  
     processor_AB AB_1_90 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_90),
       .start_in   (start_in_1_90),
       .swap_in   (swap_in_1_90),
       .op_in      (op_in_1_90),
       .pivot_in   (pivot_in_1_90),
       .start_out  (start_out_1_90),
       .swap_out   (swap_out_1_90),
       .data_out   (data_out_1_90),
       .op_out     (op_out_1_90),
       .pivot_out  (pivot_out_1_90),
       .r          (r_1_90)
     );

  // row 1, col 91

     reg start_in_1_91;
     wire start_out_1_91;

     reg swap_in_1_91;
     wire swap_out_1_91;

     reg [1:0] op_in_1_91;
     wire [1:0] op_out_1_91;

     wire r_1_91;

     reg data_in_1_91;
     wire data_out_1_91;

     reg pivot_in_1_91;
     wire pivot_out_1_91;

     always @(posedge clk) begin
         op_in_1_91 <= op_out_1_90;
         pivot_in_1_91 <= pivot_out_1_90;
         start_in_1_91 <= start_out_1_90;
         swap_in_1_91 <= swap_out_1_90;
     end

     always @(posedge clk) begin
         data_in_1_91 <= data_out_0_91;
     end
  
     processor_AB AB_1_91 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_91),
       .start_in   (start_in_1_91),
       .swap_in   (swap_in_1_91),
       .op_in      (op_in_1_91),
       .pivot_in   (pivot_in_1_91),
       .start_out  (start_out_1_91),
       .swap_out   (swap_out_1_91),
       .data_out   (data_out_1_91),
       .op_out     (op_out_1_91),
       .pivot_out  (pivot_out_1_91),
       .r          (r_1_91)
     );

  // row 1, col 92

     reg start_in_1_92;
     wire start_out_1_92;

     reg swap_in_1_92;
     wire swap_out_1_92;

     reg [1:0] op_in_1_92;
     wire [1:0] op_out_1_92;

     wire r_1_92;

     reg data_in_1_92;
     wire data_out_1_92;

     reg pivot_in_1_92;
     wire pivot_out_1_92;

     always @(posedge clk) begin
         op_in_1_92 <= op_out_1_91;
         pivot_in_1_92 <= pivot_out_1_91;
         start_in_1_92 <= start_out_1_91;
         swap_in_1_92 <= swap_out_1_91;
     end

     always @(posedge clk) begin
         data_in_1_92 <= data_out_0_92;
     end
  
     processor_AB AB_1_92 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_92),
       .start_in   (start_in_1_92),
       .swap_in   (swap_in_1_92),
       .op_in      (op_in_1_92),
       .pivot_in   (pivot_in_1_92),
       .start_out  (start_out_1_92),
       .swap_out   (swap_out_1_92),
       .data_out   (data_out_1_92),
       .op_out     (op_out_1_92),
       .pivot_out  (pivot_out_1_92),
       .r          (r_1_92)
     );

  // row 1, col 93

     reg start_in_1_93;
     wire start_out_1_93;

     reg swap_in_1_93;
     wire swap_out_1_93;

     reg [1:0] op_in_1_93;
     wire [1:0] op_out_1_93;

     wire r_1_93;

     reg data_in_1_93;
     wire data_out_1_93;

     reg pivot_in_1_93;
     wire pivot_out_1_93;

     always @(posedge clk) begin
         op_in_1_93 <= op_out_1_92;
         pivot_in_1_93 <= pivot_out_1_92;
         start_in_1_93 <= start_out_1_92;
         swap_in_1_93 <= swap_out_1_92;
     end

     always @(posedge clk) begin
         data_in_1_93 <= data_out_0_93;
     end
  
     processor_AB AB_1_93 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_93),
       .start_in   (start_in_1_93),
       .swap_in   (swap_in_1_93),
       .op_in      (op_in_1_93),
       .pivot_in   (pivot_in_1_93),
       .start_out  (start_out_1_93),
       .swap_out   (swap_out_1_93),
       .data_out   (data_out_1_93),
       .op_out     (op_out_1_93),
       .pivot_out  (pivot_out_1_93),
       .r          (r_1_93)
     );

  // row 1, col 94

     reg start_in_1_94;
     wire start_out_1_94;

     reg swap_in_1_94;
     wire swap_out_1_94;

     reg [1:0] op_in_1_94;
     wire [1:0] op_out_1_94;

     wire r_1_94;

     reg data_in_1_94;
     wire data_out_1_94;

     reg pivot_in_1_94;
     wire pivot_out_1_94;

     always @(posedge clk) begin
         op_in_1_94 <= op_out_1_93;
         pivot_in_1_94 <= pivot_out_1_93;
         start_in_1_94 <= start_out_1_93;
         swap_in_1_94 <= swap_out_1_93;
     end

     always @(posedge clk) begin
         data_in_1_94 <= data_out_0_94;
     end
  
     processor_AB AB_1_94 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_94),
       .start_in   (start_in_1_94),
       .swap_in   (swap_in_1_94),
       .op_in      (op_in_1_94),
       .pivot_in   (pivot_in_1_94),
       .start_out  (start_out_1_94),
       .swap_out   (swap_out_1_94),
       .data_out   (data_out_1_94),
       .op_out     (op_out_1_94),
       .pivot_out  (pivot_out_1_94),
       .r          (r_1_94)
     );

  // row 1, col 95

     reg start_in_1_95;
     wire start_out_1_95;

     reg swap_in_1_95;
     wire swap_out_1_95;

     reg [1:0] op_in_1_95;
     wire [1:0] op_out_1_95;

     wire r_1_95;

     reg data_in_1_95;
     wire data_out_1_95;

     reg pivot_in_1_95;
     wire pivot_out_1_95;

     always @(posedge clk) begin
         op_in_1_95 <= op_out_1_94;
         pivot_in_1_95 <= pivot_out_1_94;
         start_in_1_95 <= start_out_1_94;
         swap_in_1_95 <= swap_out_1_94;
     end

     always @(posedge clk) begin
         data_in_1_95 <= data_out_0_95;
     end
  
     processor_AB AB_1_95 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_95),
       .start_in   (start_in_1_95),
       .swap_in   (swap_in_1_95),
       .op_in      (op_in_1_95),
       .pivot_in   (pivot_in_1_95),
       .start_out  (start_out_1_95),
       .swap_out   (swap_out_1_95),
       .data_out   (data_out_1_95),
       .op_out     (op_out_1_95),
       .pivot_out  (pivot_out_1_95),
       .r          (r_1_95)
     );

  // row 1, col 96

     reg start_in_1_96;
     wire start_out_1_96;

     reg swap_in_1_96;
     wire swap_out_1_96;

     reg [1:0] op_in_1_96;
     wire [1:0] op_out_1_96;

     wire r_1_96;

     reg data_in_1_96;
     wire data_out_1_96;

     reg pivot_in_1_96;
     wire pivot_out_1_96;

     always @(posedge clk) begin
         op_in_1_96 <= op_out_1_95;
         pivot_in_1_96 <= pivot_out_1_95;
         start_in_1_96 <= start_out_1_95;
         swap_in_1_96 <= swap_out_1_95;
     end

     always @(posedge clk) begin
         data_in_1_96 <= data_out_0_96;
     end
  
     processor_AB AB_1_96 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_96),
       .start_in   (start_in_1_96),
       .swap_in   (swap_in_1_96),
       .op_in      (op_in_1_96),
       .pivot_in   (pivot_in_1_96),
       .start_out  (start_out_1_96),
       .swap_out   (swap_out_1_96),
       .data_out   (data_out_1_96),
       .op_out     (op_out_1_96),
       .pivot_out  (pivot_out_1_96),
       .r          (r_1_96)
     );

  // row 1, col 97

     reg start_in_1_97;
     wire start_out_1_97;

     reg swap_in_1_97;
     wire swap_out_1_97;

     reg [1:0] op_in_1_97;
     wire [1:0] op_out_1_97;

     wire r_1_97;

     reg data_in_1_97;
     wire data_out_1_97;

     reg pivot_in_1_97;
     wire pivot_out_1_97;

     always @(posedge clk) begin
         op_in_1_97 <= op_out_1_96;
         pivot_in_1_97 <= pivot_out_1_96;
         start_in_1_97 <= start_out_1_96;
         swap_in_1_97 <= swap_out_1_96;
     end

     always @(posedge clk) begin
         data_in_1_97 <= data_out_0_97;
     end
  
     processor_AB AB_1_97 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_97),
       .start_in   (start_in_1_97),
       .swap_in   (swap_in_1_97),
       .op_in      (op_in_1_97),
       .pivot_in   (pivot_in_1_97),
       .start_out  (start_out_1_97),
       .swap_out   (swap_out_1_97),
       .data_out   (data_out_1_97),
       .op_out     (op_out_1_97),
       .pivot_out  (pivot_out_1_97),
       .r          (r_1_97)
     );

  // row 1, col 98

     reg start_in_1_98;
     wire start_out_1_98;

     reg swap_in_1_98;
     wire swap_out_1_98;

     reg [1:0] op_in_1_98;
     wire [1:0] op_out_1_98;

     wire r_1_98;

     reg data_in_1_98;
     wire data_out_1_98;

     reg pivot_in_1_98;
     wire pivot_out_1_98;

     always @(posedge clk) begin
         op_in_1_98 <= op_out_1_97;
         pivot_in_1_98 <= pivot_out_1_97;
         start_in_1_98 <= start_out_1_97;
         swap_in_1_98 <= swap_out_1_97;
     end

     always @(posedge clk) begin
         data_in_1_98 <= data_out_0_98;
     end
  
     processor_AB AB_1_98 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_98),
       .start_in   (start_in_1_98),
       .swap_in   (swap_in_1_98),
       .op_in      (op_in_1_98),
       .pivot_in   (pivot_in_1_98),
       .start_out  (start_out_1_98),
       .swap_out   (swap_out_1_98),
       .data_out   (data_out_1_98),
       .op_out     (op_out_1_98),
       .pivot_out  (pivot_out_1_98),
       .r          (r_1_98)
     );

  // row 1, col 99

     reg start_in_1_99;
     wire start_out_1_99;

     reg swap_in_1_99;
     wire swap_out_1_99;

     reg [1:0] op_in_1_99;
     wire [1:0] op_out_1_99;

     wire r_1_99;

     reg data_in_1_99;
     wire data_out_1_99;

     reg pivot_in_1_99;
     wire pivot_out_1_99;

     always @(posedge clk) begin
         op_in_1_99 <= op_out_1_98;
         pivot_in_1_99 <= pivot_out_1_98;
         start_in_1_99 <= start_out_1_98;
         swap_in_1_99 <= swap_out_1_98;
     end

     always @(posedge clk) begin
         data_in_1_99 <= data_out_0_99;
     end
  
     processor_AB AB_1_99 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_99),
       .start_in   (start_in_1_99),
       .swap_in   (swap_in_1_99),
       .op_in      (op_in_1_99),
       .pivot_in   (pivot_in_1_99),
       .start_out  (start_out_1_99),
       .swap_out   (swap_out_1_99),
       .data_out   (data_out_1_99),
       .op_out     (op_out_1_99),
       .pivot_out  (pivot_out_1_99),
       .r          (r_1_99)
     );

  // row 1, col 100

     reg start_in_1_100;
     wire start_out_1_100;

     reg swap_in_1_100;
     wire swap_out_1_100;

     reg [1:0] op_in_1_100;
     wire [1:0] op_out_1_100;

     wire r_1_100;

     reg data_in_1_100;
     wire data_out_1_100;

     reg pivot_in_1_100;
     wire pivot_out_1_100;

     always @(posedge clk) begin
         op_in_1_100 <= op_out_1_99;
         pivot_in_1_100 <= pivot_out_1_99;
         start_in_1_100 <= start_out_1_99;
         swap_in_1_100 <= swap_out_1_99;
     end

     always @(posedge clk) begin
         data_in_1_100 <= data_out_0_100;
     end
  
     processor_AB AB_1_100 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_100),
       .start_in   (start_in_1_100),
       .swap_in   (swap_in_1_100),
       .op_in      (op_in_1_100),
       .pivot_in   (pivot_in_1_100),
       .start_out  (start_out_1_100),
       .swap_out   (swap_out_1_100),
       .data_out   (data_out_1_100),
       .op_out     (op_out_1_100),
       .pivot_out  (pivot_out_1_100),
       .r          (r_1_100)
     );

  // row 1, col 101

     reg start_in_1_101;
     wire start_out_1_101;

     reg swap_in_1_101;
     wire swap_out_1_101;

     reg [1:0] op_in_1_101;
     wire [1:0] op_out_1_101;

     wire r_1_101;

     reg data_in_1_101;
     wire data_out_1_101;

     reg pivot_in_1_101;
     wire pivot_out_1_101;

     always @(posedge clk) begin
         op_in_1_101 <= op_out_1_100;
         pivot_in_1_101 <= pivot_out_1_100;
         start_in_1_101 <= start_out_1_100;
         swap_in_1_101 <= swap_out_1_100;
     end

     always @(posedge clk) begin
         data_in_1_101 <= data_out_0_101;
     end
  
     processor_AB AB_1_101 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_101),
       .start_in   (start_in_1_101),
       .swap_in   (swap_in_1_101),
       .op_in      (op_in_1_101),
       .pivot_in   (pivot_in_1_101),
       .start_out  (start_out_1_101),
       .swap_out   (swap_out_1_101),
       .data_out   (data_out_1_101),
       .op_out     (op_out_1_101),
       .pivot_out  (pivot_out_1_101),
       .r          (r_1_101)
     );

  // row 1, col 102

     reg start_in_1_102;
     wire start_out_1_102;

     reg swap_in_1_102;
     wire swap_out_1_102;

     reg [1:0] op_in_1_102;
     wire [1:0] op_out_1_102;

     wire r_1_102;

     reg data_in_1_102;
     wire data_out_1_102;

     reg pivot_in_1_102;
     wire pivot_out_1_102;

     always @(posedge clk) begin
         op_in_1_102 <= op_out_1_101;
         pivot_in_1_102 <= pivot_out_1_101;
         start_in_1_102 <= start_out_1_101;
         swap_in_1_102 <= swap_out_1_101;
     end

     always @(posedge clk) begin
         data_in_1_102 <= data_out_0_102;
     end
  
     processor_AB AB_1_102 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_102),
       .start_in   (start_in_1_102),
       .swap_in   (swap_in_1_102),
       .op_in      (op_in_1_102),
       .pivot_in   (pivot_in_1_102),
       .start_out  (start_out_1_102),
       .swap_out   (swap_out_1_102),
       .data_out   (data_out_1_102),
       .op_out     (op_out_1_102),
       .pivot_out  (pivot_out_1_102),
       .r          (r_1_102)
     );

  // row 1, col 103

     reg start_in_1_103;
     wire start_out_1_103;

     reg swap_in_1_103;
     wire swap_out_1_103;

     reg [1:0] op_in_1_103;
     wire [1:0] op_out_1_103;

     wire r_1_103;

     reg data_in_1_103;
     wire data_out_1_103;

     reg pivot_in_1_103;
     wire pivot_out_1_103;

     always @(posedge clk) begin
         op_in_1_103 <= op_out_1_102;
         pivot_in_1_103 <= pivot_out_1_102;
         start_in_1_103 <= start_out_1_102;
         swap_in_1_103 <= swap_out_1_102;
     end

     always @(posedge clk) begin
         data_in_1_103 <= data_out_0_103;
     end
  
     processor_AB AB_1_103 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_103),
       .start_in   (start_in_1_103),
       .swap_in   (swap_in_1_103),
       .op_in      (op_in_1_103),
       .pivot_in   (pivot_in_1_103),
       .start_out  (start_out_1_103),
       .swap_out   (swap_out_1_103),
       .data_out   (data_out_1_103),
       .op_out     (op_out_1_103),
       .pivot_out  (pivot_out_1_103),
       .r          (r_1_103)
     );

  // row 1, col 104

     reg start_in_1_104;
     wire start_out_1_104;

     reg swap_in_1_104;
     wire swap_out_1_104;

     reg [1:0] op_in_1_104;
     wire [1:0] op_out_1_104;

     wire r_1_104;

     reg data_in_1_104;
     wire data_out_1_104;

     reg pivot_in_1_104;
     wire pivot_out_1_104;

     always @(posedge clk) begin
         op_in_1_104 <= op_out_1_103;
         pivot_in_1_104 <= pivot_out_1_103;
         start_in_1_104 <= start_out_1_103;
         swap_in_1_104 <= swap_out_1_103;
     end

     always @(posedge clk) begin
         data_in_1_104 <= data_out_0_104;
     end
  
     processor_AB AB_1_104 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_104),
       .start_in   (start_in_1_104),
       .swap_in   (swap_in_1_104),
       .op_in      (op_in_1_104),
       .pivot_in   (pivot_in_1_104),
       .start_out  (start_out_1_104),
       .swap_out   (swap_out_1_104),
       .data_out   (data_out_1_104),
       .op_out     (op_out_1_104),
       .pivot_out  (pivot_out_1_104),
       .r          (r_1_104)
     );

  // row 1, col 105

     reg start_in_1_105;
     wire start_out_1_105;

     reg swap_in_1_105;
     wire swap_out_1_105;

     reg [1:0] op_in_1_105;
     wire [1:0] op_out_1_105;

     wire r_1_105;

     reg data_in_1_105;
     wire data_out_1_105;

     reg pivot_in_1_105;
     wire pivot_out_1_105;

     always @(posedge clk) begin
         op_in_1_105 <= op_out_1_104;
         pivot_in_1_105 <= pivot_out_1_104;
         start_in_1_105 <= start_out_1_104;
         swap_in_1_105 <= swap_out_1_104;
     end

     always @(posedge clk) begin
         data_in_1_105 <= data_out_0_105;
     end
  
     processor_AB AB_1_105 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_105),
       .start_in   (start_in_1_105),
       .swap_in   (swap_in_1_105),
       .op_in      (op_in_1_105),
       .pivot_in   (pivot_in_1_105),
       .start_out  (start_out_1_105),
       .swap_out   (swap_out_1_105),
       .data_out   (data_out_1_105),
       .op_out     (op_out_1_105),
       .pivot_out  (pivot_out_1_105),
       .r          (r_1_105)
     );

  // row 1, col 106

     reg start_in_1_106;
     wire start_out_1_106;

     reg swap_in_1_106;
     wire swap_out_1_106;

     reg [1:0] op_in_1_106;
     wire [1:0] op_out_1_106;

     wire r_1_106;

     reg data_in_1_106;
     wire data_out_1_106;

     reg pivot_in_1_106;
     wire pivot_out_1_106;

     always @(posedge clk) begin
         op_in_1_106 <= op_out_1_105;
         pivot_in_1_106 <= pivot_out_1_105;
         start_in_1_106 <= start_out_1_105;
         swap_in_1_106 <= swap_out_1_105;
     end

     always @(posedge clk) begin
         data_in_1_106 <= data_out_0_106;
     end
  
     processor_AB AB_1_106 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_106),
       .start_in   (start_in_1_106),
       .swap_in   (swap_in_1_106),
       .op_in      (op_in_1_106),
       .pivot_in   (pivot_in_1_106),
       .start_out  (start_out_1_106),
       .swap_out   (swap_out_1_106),
       .data_out   (data_out_1_106),
       .op_out     (op_out_1_106),
       .pivot_out  (pivot_out_1_106),
       .r          (r_1_106)
     );

  // row 1, col 107

     reg start_in_1_107;
     wire start_out_1_107;

     reg swap_in_1_107;
     wire swap_out_1_107;

     reg [1:0] op_in_1_107;
     wire [1:0] op_out_1_107;

     wire r_1_107;

     reg data_in_1_107;
     wire data_out_1_107;

     reg pivot_in_1_107;
     wire pivot_out_1_107;

     always @(posedge clk) begin
         op_in_1_107 <= op_out_1_106;
         pivot_in_1_107 <= pivot_out_1_106;
         start_in_1_107 <= start_out_1_106;
         swap_in_1_107 <= swap_out_1_106;
     end

     always @(posedge clk) begin
         data_in_1_107 <= data_out_0_107;
     end
  
     processor_AB AB_1_107 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_107),
       .start_in   (start_in_1_107),
       .swap_in   (swap_in_1_107),
       .op_in      (op_in_1_107),
       .pivot_in   (pivot_in_1_107),
       .start_out  (start_out_1_107),
       .swap_out   (swap_out_1_107),
       .data_out   (data_out_1_107),
       .op_out     (op_out_1_107),
       .pivot_out  (pivot_out_1_107),
       .r          (r_1_107)
     );

  // row 1, col 108

     reg start_in_1_108;
     wire start_out_1_108;

     reg swap_in_1_108;
     wire swap_out_1_108;

     reg [1:0] op_in_1_108;
     wire [1:0] op_out_1_108;

     wire r_1_108;

     reg data_in_1_108;
     wire data_out_1_108;

     reg pivot_in_1_108;
     wire pivot_out_1_108;

     always @(posedge clk) begin
         op_in_1_108 <= op_out_1_107;
         pivot_in_1_108 <= pivot_out_1_107;
         start_in_1_108 <= start_out_1_107;
         swap_in_1_108 <= swap_out_1_107;
     end

     always @(posedge clk) begin
         data_in_1_108 <= data_out_0_108;
     end
  
     processor_AB AB_1_108 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_108),
       .start_in   (start_in_1_108),
       .swap_in   (swap_in_1_108),
       .op_in      (op_in_1_108),
       .pivot_in   (pivot_in_1_108),
       .start_out  (start_out_1_108),
       .swap_out   (swap_out_1_108),
       .data_out   (data_out_1_108),
       .op_out     (op_out_1_108),
       .pivot_out  (pivot_out_1_108),
       .r          (r_1_108)
     );

  // row 1, col 109

     reg start_in_1_109;
     wire start_out_1_109;

     reg swap_in_1_109;
     wire swap_out_1_109;

     reg [1:0] op_in_1_109;
     wire [1:0] op_out_1_109;

     wire r_1_109;

     reg data_in_1_109;
     wire data_out_1_109;

     reg pivot_in_1_109;
     wire pivot_out_1_109;

     always @(posedge clk) begin
         op_in_1_109 <= op_out_1_108;
         pivot_in_1_109 <= pivot_out_1_108;
         start_in_1_109 <= start_out_1_108;
         swap_in_1_109 <= swap_out_1_108;
     end

     always @(posedge clk) begin
         data_in_1_109 <= data_out_0_109;
     end
  
     processor_AB AB_1_109 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_109),
       .start_in   (start_in_1_109),
       .swap_in   (swap_in_1_109),
       .op_in      (op_in_1_109),
       .pivot_in   (pivot_in_1_109),
       .start_out  (start_out_1_109),
       .swap_out   (swap_out_1_109),
       .data_out   (data_out_1_109),
       .op_out     (op_out_1_109),
       .pivot_out  (pivot_out_1_109),
       .r          (r_1_109)
     );

  // row 1, col 110

     reg start_in_1_110;
     wire start_out_1_110;

     reg swap_in_1_110;
     wire swap_out_1_110;

     reg [1:0] op_in_1_110;
     wire [1:0] op_out_1_110;

     wire r_1_110;

     reg data_in_1_110;
     wire data_out_1_110;

     reg pivot_in_1_110;
     wire pivot_out_1_110;

     always @(posedge clk) begin
         op_in_1_110 <= op_out_1_109;
         pivot_in_1_110 <= pivot_out_1_109;
         start_in_1_110 <= start_out_1_109;
         swap_in_1_110 <= swap_out_1_109;
     end

     always @(posedge clk) begin
         data_in_1_110 <= data_out_0_110;
     end
  
     processor_AB AB_1_110 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_110),
       .start_in   (start_in_1_110),
       .swap_in   (swap_in_1_110),
       .op_in      (op_in_1_110),
       .pivot_in   (pivot_in_1_110),
       .start_out  (start_out_1_110),
       .swap_out   (swap_out_1_110),
       .data_out   (data_out_1_110),
       .op_out     (op_out_1_110),
       .pivot_out  (pivot_out_1_110),
       .r          (r_1_110)
     );

  // row 1, col 111

     reg start_in_1_111;
     wire start_out_1_111;

     reg swap_in_1_111;
     wire swap_out_1_111;

     reg [1:0] op_in_1_111;
     wire [1:0] op_out_1_111;

     wire r_1_111;

     reg data_in_1_111;
     wire data_out_1_111;

     reg pivot_in_1_111;
     wire pivot_out_1_111;

     always @(posedge clk) begin
         op_in_1_111 <= op_out_1_110;
         pivot_in_1_111 <= pivot_out_1_110;
         start_in_1_111 <= start_out_1_110;
         swap_in_1_111 <= swap_out_1_110;
     end

     always @(posedge clk) begin
         data_in_1_111 <= data_out_0_111;
     end
  
     processor_AB AB_1_111 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_111),
       .start_in   (start_in_1_111),
       .swap_in   (swap_in_1_111),
       .op_in      (op_in_1_111),
       .pivot_in   (pivot_in_1_111),
       .start_out  (start_out_1_111),
       .swap_out   (swap_out_1_111),
       .data_out   (data_out_1_111),
       .op_out     (op_out_1_111),
       .pivot_out  (pivot_out_1_111),
       .r          (r_1_111)
     );

  // row 1, col 112

     reg start_in_1_112;
     wire start_out_1_112;

     reg swap_in_1_112;
     wire swap_out_1_112;

     reg [1:0] op_in_1_112;
     wire [1:0] op_out_1_112;

     wire r_1_112;

     reg data_in_1_112;
     wire data_out_1_112;

     reg pivot_in_1_112;
     wire pivot_out_1_112;

     always @(posedge clk) begin
         op_in_1_112 <= op_out_1_111;
         pivot_in_1_112 <= pivot_out_1_111;
         start_in_1_112 <= start_out_1_111;
         swap_in_1_112 <= swap_out_1_111;
     end

     always @(posedge clk) begin
         data_in_1_112 <= data_out_0_112;
     end
  
     processor_AB AB_1_112 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_112),
       .start_in   (start_in_1_112),
       .swap_in   (swap_in_1_112),
       .op_in      (op_in_1_112),
       .pivot_in   (pivot_in_1_112),
       .start_out  (start_out_1_112),
       .swap_out   (swap_out_1_112),
       .data_out   (data_out_1_112),
       .op_out     (op_out_1_112),
       .pivot_out  (pivot_out_1_112),
       .r          (r_1_112)
     );

  // row 1, col 113

     reg start_in_1_113;
     wire start_out_1_113;

     reg swap_in_1_113;
     wire swap_out_1_113;

     reg [1:0] op_in_1_113;
     wire [1:0] op_out_1_113;

     wire r_1_113;

     reg data_in_1_113;
     wire data_out_1_113;

     reg pivot_in_1_113;
     wire pivot_out_1_113;

     always @(posedge clk) begin
         op_in_1_113 <= op_out_1_112;
         pivot_in_1_113 <= pivot_out_1_112;
         start_in_1_113 <= start_out_1_112;
         swap_in_1_113 <= swap_out_1_112;
     end

     always @(posedge clk) begin
         data_in_1_113 <= data_out_0_113;
     end
  
     processor_AB AB_1_113 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_113),
       .start_in   (start_in_1_113),
       .swap_in   (swap_in_1_113),
       .op_in      (op_in_1_113),
       .pivot_in   (pivot_in_1_113),
       .start_out  (start_out_1_113),
       .swap_out   (swap_out_1_113),
       .data_out   (data_out_1_113),
       .op_out     (op_out_1_113),
       .pivot_out  (pivot_out_1_113),
       .r          (r_1_113)
     );

  // row 1, col 114

     reg start_in_1_114;
     wire start_out_1_114;

     reg swap_in_1_114;
     wire swap_out_1_114;

     reg [1:0] op_in_1_114;
     wire [1:0] op_out_1_114;

     wire r_1_114;

     reg data_in_1_114;
     wire data_out_1_114;

     reg pivot_in_1_114;
     wire pivot_out_1_114;

     always @(posedge clk) begin
         op_in_1_114 <= op_out_1_113;
         pivot_in_1_114 <= pivot_out_1_113;
         start_in_1_114 <= start_out_1_113;
         swap_in_1_114 <= swap_out_1_113;
     end

     always @(posedge clk) begin
         data_in_1_114 <= data_out_0_114;
     end
  
     processor_AB AB_1_114 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_114),
       .start_in   (start_in_1_114),
       .swap_in   (swap_in_1_114),
       .op_in      (op_in_1_114),
       .pivot_in   (pivot_in_1_114),
       .start_out  (start_out_1_114),
       .swap_out   (swap_out_1_114),
       .data_out   (data_out_1_114),
       .op_out     (op_out_1_114),
       .pivot_out  (pivot_out_1_114),
       .r          (r_1_114)
     );

  // row 1, col 115

     reg start_in_1_115;
     wire start_out_1_115;

     reg swap_in_1_115;
     wire swap_out_1_115;

     reg [1:0] op_in_1_115;
     wire [1:0] op_out_1_115;

     wire r_1_115;

     reg data_in_1_115;
     wire data_out_1_115;

     reg pivot_in_1_115;
     wire pivot_out_1_115;

     always @(posedge clk) begin
         op_in_1_115 <= op_out_1_114;
         pivot_in_1_115 <= pivot_out_1_114;
         start_in_1_115 <= start_out_1_114;
         swap_in_1_115 <= swap_out_1_114;
     end

     always @(posedge clk) begin
         data_in_1_115 <= data_out_0_115;
     end
  
     processor_AB AB_1_115 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_115),
       .start_in   (start_in_1_115),
       .swap_in   (swap_in_1_115),
       .op_in      (op_in_1_115),
       .pivot_in   (pivot_in_1_115),
       .start_out  (start_out_1_115),
       .swap_out   (swap_out_1_115),
       .data_out   (data_out_1_115),
       .op_out     (op_out_1_115),
       .pivot_out  (pivot_out_1_115),
       .r          (r_1_115)
     );

  // row 1, col 116

     reg start_in_1_116;
     wire start_out_1_116;

     reg swap_in_1_116;
     wire swap_out_1_116;

     reg [1:0] op_in_1_116;
     wire [1:0] op_out_1_116;

     wire r_1_116;

     reg data_in_1_116;
     wire data_out_1_116;

     reg pivot_in_1_116;
     wire pivot_out_1_116;

     always @(posedge clk) begin
         op_in_1_116 <= op_out_1_115;
         pivot_in_1_116 <= pivot_out_1_115;
         start_in_1_116 <= start_out_1_115;
         swap_in_1_116 <= swap_out_1_115;
     end

     always @(posedge clk) begin
         data_in_1_116 <= data_out_0_116;
     end
  
     processor_AB AB_1_116 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_116),
       .start_in   (start_in_1_116),
       .swap_in   (swap_in_1_116),
       .op_in      (op_in_1_116),
       .pivot_in   (pivot_in_1_116),
       .start_out  (start_out_1_116),
       .swap_out   (swap_out_1_116),
       .data_out   (data_out_1_116),
       .op_out     (op_out_1_116),
       .pivot_out  (pivot_out_1_116),
       .r          (r_1_116)
     );

  // row 1, col 117

     reg start_in_1_117;
     wire start_out_1_117;

     reg swap_in_1_117;
     wire swap_out_1_117;

     reg [1:0] op_in_1_117;
     wire [1:0] op_out_1_117;

     wire r_1_117;

     reg data_in_1_117;
     wire data_out_1_117;

     reg pivot_in_1_117;
     wire pivot_out_1_117;

     always @(posedge clk) begin
         op_in_1_117 <= op_out_1_116;
         pivot_in_1_117 <= pivot_out_1_116;
         start_in_1_117 <= start_out_1_116;
         swap_in_1_117 <= swap_out_1_116;
     end

     always @(posedge clk) begin
         data_in_1_117 <= data_out_0_117;
     end
  
     processor_AB AB_1_117 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_117),
       .start_in   (start_in_1_117),
       .swap_in   (swap_in_1_117),
       .op_in      (op_in_1_117),
       .pivot_in   (pivot_in_1_117),
       .start_out  (start_out_1_117),
       .swap_out   (swap_out_1_117),
       .data_out   (data_out_1_117),
       .op_out     (op_out_1_117),
       .pivot_out  (pivot_out_1_117),
       .r          (r_1_117)
     );

  // row 1, col 118

     reg start_in_1_118;
     wire start_out_1_118;

     reg swap_in_1_118;
     wire swap_out_1_118;

     reg [1:0] op_in_1_118;
     wire [1:0] op_out_1_118;

     wire r_1_118;

     reg data_in_1_118;
     wire data_out_1_118;

     reg pivot_in_1_118;
     wire pivot_out_1_118;

     always @(posedge clk) begin
         op_in_1_118 <= op_out_1_117;
         pivot_in_1_118 <= pivot_out_1_117;
         start_in_1_118 <= start_out_1_117;
         swap_in_1_118 <= swap_out_1_117;
     end

     always @(posedge clk) begin
         data_in_1_118 <= data_out_0_118;
     end
  
     processor_AB AB_1_118 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_118),
       .start_in   (start_in_1_118),
       .swap_in   (swap_in_1_118),
       .op_in      (op_in_1_118),
       .pivot_in   (pivot_in_1_118),
       .start_out  (start_out_1_118),
       .swap_out   (swap_out_1_118),
       .data_out   (data_out_1_118),
       .op_out     (op_out_1_118),
       .pivot_out  (pivot_out_1_118),
       .r          (r_1_118)
     );

  // row 1, col 119

     reg start_in_1_119;
     wire start_out_1_119;

     reg swap_in_1_119;
     wire swap_out_1_119;

     reg [1:0] op_in_1_119;
     wire [1:0] op_out_1_119;

     wire r_1_119;

     reg data_in_1_119;
     wire data_out_1_119;

     reg pivot_in_1_119;
     wire pivot_out_1_119;

     always @(posedge clk) begin
         op_in_1_119 <= op_out_1_118;
         pivot_in_1_119 <= pivot_out_1_118;
         start_in_1_119 <= start_out_1_118;
         swap_in_1_119 <= swap_out_1_118;
     end

     always @(posedge clk) begin
         data_in_1_119 <= data_out_0_119;
     end
  
     processor_AB AB_1_119 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_119),
       .start_in   (start_in_1_119),
       .swap_in   (swap_in_1_119),
       .op_in      (op_in_1_119),
       .pivot_in   (pivot_in_1_119),
       .start_out  (start_out_1_119),
       .swap_out   (swap_out_1_119),
       .data_out   (data_out_1_119),
       .op_out     (op_out_1_119),
       .pivot_out  (pivot_out_1_119),
       .r          (r_1_119)
     );

  // row 1, col 120

     reg start_in_1_120;
     wire start_out_1_120;

     reg swap_in_1_120;
     wire swap_out_1_120;

     reg [1:0] op_in_1_120;
     wire [1:0] op_out_1_120;

     wire r_1_120;

     reg data_in_1_120;
     wire data_out_1_120;

     reg pivot_in_1_120;
     wire pivot_out_1_120;

     always @(posedge clk) begin
         op_in_1_120 <= op_out_1_119;
         pivot_in_1_120 <= pivot_out_1_119;
         start_in_1_120 <= start_out_1_119;
         swap_in_1_120 <= swap_out_1_119;
     end

     always @(posedge clk) begin
         data_in_1_120 <= data_out_0_120;
     end
  
     processor_AB AB_1_120 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_120),
       .start_in   (start_in_1_120),
       .swap_in   (swap_in_1_120),
       .op_in      (op_in_1_120),
       .pivot_in   (pivot_in_1_120),
       .start_out  (start_out_1_120),
       .swap_out   (swap_out_1_120),
       .data_out   (data_out_1_120),
       .op_out     (op_out_1_120),
       .pivot_out  (pivot_out_1_120),
       .r          (r_1_120)
     );

  // row 1, col 121

     reg start_in_1_121;
     wire start_out_1_121;

     reg swap_in_1_121;
     wire swap_out_1_121;

     reg [1:0] op_in_1_121;
     wire [1:0] op_out_1_121;

     wire r_1_121;

     reg data_in_1_121;
     wire data_out_1_121;

     reg pivot_in_1_121;
     wire pivot_out_1_121;

     always @(posedge clk) begin
         op_in_1_121 <= op_out_1_120;
         pivot_in_1_121 <= pivot_out_1_120;
         start_in_1_121 <= start_out_1_120;
         swap_in_1_121 <= swap_out_1_120;
     end

     always @(posedge clk) begin
         data_in_1_121 <= data_out_0_121;
     end
  
     processor_AB AB_1_121 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_121),
       .start_in   (start_in_1_121),
       .swap_in   (swap_in_1_121),
       .op_in      (op_in_1_121),
       .pivot_in   (pivot_in_1_121),
       .start_out  (start_out_1_121),
       .swap_out   (swap_out_1_121),
       .data_out   (data_out_1_121),
       .op_out     (op_out_1_121),
       .pivot_out  (pivot_out_1_121),
       .r          (r_1_121)
     );

  // row 1, col 122

     reg start_in_1_122;
     wire start_out_1_122;

     reg swap_in_1_122;
     wire swap_out_1_122;

     reg [1:0] op_in_1_122;
     wire [1:0] op_out_1_122;

     wire r_1_122;

     reg data_in_1_122;
     wire data_out_1_122;

     reg pivot_in_1_122;
     wire pivot_out_1_122;

     always @(posedge clk) begin
         op_in_1_122 <= op_out_1_121;
         pivot_in_1_122 <= pivot_out_1_121;
         start_in_1_122 <= start_out_1_121;
         swap_in_1_122 <= swap_out_1_121;
     end

     always @(posedge clk) begin
         data_in_1_122 <= data_out_0_122;
     end
  
     processor_AB AB_1_122 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_122),
       .start_in   (start_in_1_122),
       .swap_in   (swap_in_1_122),
       .op_in      (op_in_1_122),
       .pivot_in   (pivot_in_1_122),
       .start_out  (start_out_1_122),
       .swap_out   (swap_out_1_122),
       .data_out   (data_out_1_122),
       .op_out     (op_out_1_122),
       .pivot_out  (pivot_out_1_122),
       .r          (r_1_122)
     );

  // row 1, col 123

     reg start_in_1_123;
     wire start_out_1_123;

     reg swap_in_1_123;
     wire swap_out_1_123;

     reg [1:0] op_in_1_123;
     wire [1:0] op_out_1_123;

     wire r_1_123;

     reg data_in_1_123;
     wire data_out_1_123;

     reg pivot_in_1_123;
     wire pivot_out_1_123;

     always @(posedge clk) begin
         op_in_1_123 <= op_out_1_122;
         pivot_in_1_123 <= pivot_out_1_122;
         start_in_1_123 <= start_out_1_122;
         swap_in_1_123 <= swap_out_1_122;
     end

     always @(posedge clk) begin
         data_in_1_123 <= data_out_0_123;
     end
  
     processor_AB AB_1_123 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_123),
       .start_in   (start_in_1_123),
       .swap_in   (swap_in_1_123),
       .op_in      (op_in_1_123),
       .pivot_in   (pivot_in_1_123),
       .start_out  (start_out_1_123),
       .swap_out   (swap_out_1_123),
       .data_out   (data_out_1_123),
       .op_out     (op_out_1_123),
       .pivot_out  (pivot_out_1_123),
       .r          (r_1_123)
     );

  // row 1, col 124

     reg start_in_1_124;
     wire start_out_1_124;

     reg swap_in_1_124;
     wire swap_out_1_124;

     reg [1:0] op_in_1_124;
     wire [1:0] op_out_1_124;

     wire r_1_124;

     reg data_in_1_124;
     wire data_out_1_124;

     reg pivot_in_1_124;
     wire pivot_out_1_124;

     always @(posedge clk) begin
         op_in_1_124 <= op_out_1_123;
         pivot_in_1_124 <= pivot_out_1_123;
         start_in_1_124 <= start_out_1_123;
         swap_in_1_124 <= swap_out_1_123;
     end

     always @(posedge clk) begin
         data_in_1_124 <= data_out_0_124;
     end
  
     processor_AB AB_1_124 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_124),
       .start_in   (start_in_1_124),
       .swap_in   (swap_in_1_124),
       .op_in      (op_in_1_124),
       .pivot_in   (pivot_in_1_124),
       .start_out  (start_out_1_124),
       .swap_out   (swap_out_1_124),
       .data_out   (data_out_1_124),
       .op_out     (op_out_1_124),
       .pivot_out  (pivot_out_1_124),
       .r          (r_1_124)
     );

  // row 1, col 125

     reg start_in_1_125;
     wire start_out_1_125;

     reg swap_in_1_125;
     wire swap_out_1_125;

     reg [1:0] op_in_1_125;
     wire [1:0] op_out_1_125;

     wire r_1_125;

     reg data_in_1_125;
     wire data_out_1_125;

     reg pivot_in_1_125;
     wire pivot_out_1_125;

     always @(posedge clk) begin
         op_in_1_125 <= op_out_1_124;
         pivot_in_1_125 <= pivot_out_1_124;
         start_in_1_125 <= start_out_1_124;
         swap_in_1_125 <= swap_out_1_124;
     end

     always @(posedge clk) begin
         data_in_1_125 <= data_out_0_125;
     end
  
     processor_AB AB_1_125 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_125),
       .start_in   (start_in_1_125),
       .swap_in   (swap_in_1_125),
       .op_in      (op_in_1_125),
       .pivot_in   (pivot_in_1_125),
       .start_out  (start_out_1_125),
       .swap_out   (swap_out_1_125),
       .data_out   (data_out_1_125),
       .op_out     (op_out_1_125),
       .pivot_out  (pivot_out_1_125),
       .r          (r_1_125)
     );

  // row 1, col 126

     reg start_in_1_126;
     wire start_out_1_126;

     reg swap_in_1_126;
     wire swap_out_1_126;

     reg [1:0] op_in_1_126;
     wire [1:0] op_out_1_126;

     wire r_1_126;

     reg data_in_1_126;
     wire data_out_1_126;

     reg pivot_in_1_126;
     wire pivot_out_1_126;

     always @(posedge clk) begin
         op_in_1_126 <= op_out_1_125;
         pivot_in_1_126 <= pivot_out_1_125;
         start_in_1_126 <= start_out_1_125;
         swap_in_1_126 <= swap_out_1_125;
     end

     always @(posedge clk) begin
         data_in_1_126 <= data_out_0_126;
     end
  
     processor_AB AB_1_126 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_126),
       .start_in   (start_in_1_126),
       .swap_in   (swap_in_1_126),
       .op_in      (op_in_1_126),
       .pivot_in   (pivot_in_1_126),
       .start_out  (start_out_1_126),
       .swap_out   (swap_out_1_126),
       .data_out   (data_out_1_126),
       .op_out     (op_out_1_126),
       .pivot_out  (pivot_out_1_126),
       .r          (r_1_126)
     );

  // row 1, col 127

     reg start_in_1_127;
     wire start_out_1_127;

     reg swap_in_1_127;
     wire swap_out_1_127;

     reg [1:0] op_in_1_127;
     wire [1:0] op_out_1_127;

     wire r_1_127;

     reg data_in_1_127;
     wire data_out_1_127;

     reg pivot_in_1_127;
     wire pivot_out_1_127;

     always @(posedge clk) begin
         op_in_1_127 <= op_out_1_126;
         pivot_in_1_127 <= pivot_out_1_126;
         start_in_1_127 <= start_out_1_126;
         swap_in_1_127 <= swap_out_1_126;
     end

     always @(posedge clk) begin
         data_in_1_127 <= data_out_0_127;
     end
  
     processor_AB AB_1_127 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_127),
       .start_in   (start_in_1_127),
       .swap_in   (swap_in_1_127),
       .op_in      (op_in_1_127),
       .pivot_in   (pivot_in_1_127),
       .start_out  (start_out_1_127),
       .swap_out   (swap_out_1_127),
       .data_out   (data_out_1_127),
       .op_out     (op_out_1_127),
       .pivot_out  (pivot_out_1_127),
       .r          (r_1_127)
     );

  // row 1, col 128

     reg start_in_1_128;
     wire start_out_1_128;

     reg swap_in_1_128;
     wire swap_out_1_128;

     reg [1:0] op_in_1_128;
     wire [1:0] op_out_1_128;

     wire r_1_128;

     reg data_in_1_128;
     wire data_out_1_128;

     reg pivot_in_1_128;
     wire pivot_out_1_128;

     always @(posedge clk) begin
         op_in_1_128 <= op_out_1_127;
         pivot_in_1_128 <= pivot_out_1_127;
         start_in_1_128 <= start_out_1_127;
         swap_in_1_128 <= swap_out_1_127;
     end

     always @(posedge clk) begin
         data_in_1_128 <= data_out_0_128;
     end
  
     processor_AB AB_1_128 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_128),
       .start_in   (start_in_1_128),
       .swap_in   (swap_in_1_128),
       .op_in      (op_in_1_128),
       .pivot_in   (pivot_in_1_128),
       .start_out  (start_out_1_128),
       .swap_out   (swap_out_1_128),
       .data_out   (data_out_1_128),
       .op_out     (op_out_1_128),
       .pivot_out  (pivot_out_1_128),
       .r          (r_1_128)
     );

  // row 1, col 129

     reg start_in_1_129;
     wire start_out_1_129;

     reg swap_in_1_129;
     wire swap_out_1_129;

     reg [1:0] op_in_1_129;
     wire [1:0] op_out_1_129;

     wire r_1_129;

     reg data_in_1_129;
     wire data_out_1_129;

     reg pivot_in_1_129;
     wire pivot_out_1_129;

     always @(posedge clk) begin
         op_in_1_129 <= op_out_1_128;
         pivot_in_1_129 <= pivot_out_1_128;
         start_in_1_129 <= start_out_1_128;
         swap_in_1_129 <= swap_out_1_128;
     end

     always @(posedge clk) begin
         data_in_1_129 <= data_out_0_129;
     end
  
     processor_AB AB_1_129 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_129),
       .start_in   (start_in_1_129),
       .swap_in   (swap_in_1_129),
       .op_in      (op_in_1_129),
       .pivot_in   (pivot_in_1_129),
       .start_out  (start_out_1_129),
       .swap_out   (swap_out_1_129),
       .data_out   (data_out_1_129),
       .op_out     (op_out_1_129),
       .pivot_out  (pivot_out_1_129),
       .r          (r_1_129)
     );

  // row 1, col 130

     reg start_in_1_130;
     wire start_out_1_130;

     reg swap_in_1_130;
     wire swap_out_1_130;

     reg [1:0] op_in_1_130;
     wire [1:0] op_out_1_130;

     wire r_1_130;

     reg data_in_1_130;
     wire data_out_1_130;

     reg pivot_in_1_130;
     wire pivot_out_1_130;

     always @(posedge clk) begin
         op_in_1_130 <= op_out_1_129;
         pivot_in_1_130 <= pivot_out_1_129;
         start_in_1_130 <= start_out_1_129;
         swap_in_1_130 <= swap_out_1_129;
     end

     always @(posedge clk) begin
         data_in_1_130 <= data_out_0_130;
     end
  
     processor_AB AB_1_130 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_130),
       .start_in   (start_in_1_130),
       .swap_in   (swap_in_1_130),
       .op_in      (op_in_1_130),
       .pivot_in   (pivot_in_1_130),
       .start_out  (start_out_1_130),
       .swap_out   (swap_out_1_130),
       .data_out   (data_out_1_130),
       .op_out     (op_out_1_130),
       .pivot_out  (pivot_out_1_130),
       .r          (r_1_130)
     );

  // row 1, col 131

     reg start_in_1_131;
     wire start_out_1_131;

     reg swap_in_1_131;
     wire swap_out_1_131;

     reg [1:0] op_in_1_131;
     wire [1:0] op_out_1_131;

     wire r_1_131;

     reg data_in_1_131;
     wire data_out_1_131;

     reg pivot_in_1_131;
     wire pivot_out_1_131;

     always @(posedge clk) begin
         op_in_1_131 <= op_out_1_130;
         pivot_in_1_131 <= pivot_out_1_130;
         start_in_1_131 <= start_out_1_130;
         swap_in_1_131 <= swap_out_1_130;
     end

     always @(posedge clk) begin
         data_in_1_131 <= data_out_0_131;
     end
  
     processor_AB AB_1_131 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_131),
       .start_in   (start_in_1_131),
       .swap_in   (swap_in_1_131),
       .op_in      (op_in_1_131),
       .pivot_in   (pivot_in_1_131),
       .start_out  (start_out_1_131),
       .swap_out   (swap_out_1_131),
       .data_out   (data_out_1_131),
       .op_out     (op_out_1_131),
       .pivot_out  (pivot_out_1_131),
       .r          (r_1_131)
     );

  // row 1, col 132

     reg start_in_1_132;
     wire start_out_1_132;

     reg swap_in_1_132;
     wire swap_out_1_132;

     reg [1:0] op_in_1_132;
     wire [1:0] op_out_1_132;

     wire r_1_132;

     reg data_in_1_132;
     wire data_out_1_132;

     reg pivot_in_1_132;
     wire pivot_out_1_132;

     always @(posedge clk) begin
         op_in_1_132 <= op_out_1_131;
         pivot_in_1_132 <= pivot_out_1_131;
         start_in_1_132 <= start_out_1_131;
         swap_in_1_132 <= swap_out_1_131;
     end

     always @(posedge clk) begin
         data_in_1_132 <= data_out_0_132;
     end
  
     processor_AB AB_1_132 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_132),
       .start_in   (start_in_1_132),
       .swap_in   (swap_in_1_132),
       .op_in      (op_in_1_132),
       .pivot_in   (pivot_in_1_132),
       .start_out  (start_out_1_132),
       .swap_out   (swap_out_1_132),
       .data_out   (data_out_1_132),
       .op_out     (op_out_1_132),
       .pivot_out  (pivot_out_1_132),
       .r          (r_1_132)
     );

  // row 1, col 133

     reg start_in_1_133;
     wire start_out_1_133;

     reg swap_in_1_133;
     wire swap_out_1_133;

     reg [1:0] op_in_1_133;
     wire [1:0] op_out_1_133;

     wire r_1_133;

     reg data_in_1_133;
     wire data_out_1_133;

     reg pivot_in_1_133;
     wire pivot_out_1_133;

     always @(posedge clk) begin
         op_in_1_133 <= op_out_1_132;
         pivot_in_1_133 <= pivot_out_1_132;
         start_in_1_133 <= start_out_1_132;
         swap_in_1_133 <= swap_out_1_132;
     end

     always @(posedge clk) begin
         data_in_1_133 <= data_out_0_133;
     end
  
     processor_AB AB_1_133 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_133),
       .start_in   (start_in_1_133),
       .swap_in   (swap_in_1_133),
       .op_in      (op_in_1_133),
       .pivot_in   (pivot_in_1_133),
       .start_out  (start_out_1_133),
       .swap_out   (swap_out_1_133),
       .data_out   (data_out_1_133),
       .op_out     (op_out_1_133),
       .pivot_out  (pivot_out_1_133),
       .r          (r_1_133)
     );

  // row 1, col 134

     reg start_in_1_134;
     wire start_out_1_134;

     reg swap_in_1_134;
     wire swap_out_1_134;

     reg [1:0] op_in_1_134;
     wire [1:0] op_out_1_134;

     wire r_1_134;

     reg data_in_1_134;
     wire data_out_1_134;

     reg pivot_in_1_134;
     wire pivot_out_1_134;

     always @(posedge clk) begin
         op_in_1_134 <= op_out_1_133;
         pivot_in_1_134 <= pivot_out_1_133;
         start_in_1_134 <= start_out_1_133;
         swap_in_1_134 <= swap_out_1_133;
     end

     always @(posedge clk) begin
         data_in_1_134 <= data_out_0_134;
     end
  
     processor_AB AB_1_134 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_134),
       .start_in   (start_in_1_134),
       .swap_in   (swap_in_1_134),
       .op_in      (op_in_1_134),
       .pivot_in   (pivot_in_1_134),
       .start_out  (start_out_1_134),
       .swap_out   (swap_out_1_134),
       .data_out   (data_out_1_134),
       .op_out     (op_out_1_134),
       .pivot_out  (pivot_out_1_134),
       .r          (r_1_134)
     );

  // row 1, col 135

     reg start_in_1_135;
     wire start_out_1_135;

     reg swap_in_1_135;
     wire swap_out_1_135;

     reg [1:0] op_in_1_135;
     wire [1:0] op_out_1_135;

     wire r_1_135;

     reg data_in_1_135;
     wire data_out_1_135;

     reg pivot_in_1_135;
     wire pivot_out_1_135;

     always @(posedge clk) begin
         op_in_1_135 <= op_out_1_134;
         pivot_in_1_135 <= pivot_out_1_134;
         start_in_1_135 <= start_out_1_134;
         swap_in_1_135 <= swap_out_1_134;
     end

     always @(posedge clk) begin
         data_in_1_135 <= data_out_0_135;
     end
  
     processor_AB AB_1_135 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_135),
       .start_in   (start_in_1_135),
       .swap_in   (swap_in_1_135),
       .op_in      (op_in_1_135),
       .pivot_in   (pivot_in_1_135),
       .start_out  (start_out_1_135),
       .swap_out   (swap_out_1_135),
       .data_out   (data_out_1_135),
       .op_out     (op_out_1_135),
       .pivot_out  (pivot_out_1_135),
       .r          (r_1_135)
     );

  // row 1, col 136

     reg start_in_1_136;
     wire start_out_1_136;

     reg swap_in_1_136;
     wire swap_out_1_136;

     reg [1:0] op_in_1_136;
     wire [1:0] op_out_1_136;

     wire r_1_136;

     reg data_in_1_136;
     wire data_out_1_136;

     reg pivot_in_1_136;
     wire pivot_out_1_136;

     always @(posedge clk) begin
         op_in_1_136 <= op_out_1_135;
         pivot_in_1_136 <= pivot_out_1_135;
         start_in_1_136 <= start_out_1_135;
         swap_in_1_136 <= swap_out_1_135;
     end

     always @(posedge clk) begin
         data_in_1_136 <= data_out_0_136;
     end
  
     processor_AB AB_1_136 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_136),
       .start_in   (start_in_1_136),
       .swap_in   (swap_in_1_136),
       .op_in      (op_in_1_136),
       .pivot_in   (pivot_in_1_136),
       .start_out  (start_out_1_136),
       .swap_out   (swap_out_1_136),
       .data_out   (data_out_1_136),
       .op_out     (op_out_1_136),
       .pivot_out  (pivot_out_1_136),
       .r          (r_1_136)
     );

  // row 1, col 137

     reg start_in_1_137;
     wire start_out_1_137;

     reg swap_in_1_137;
     wire swap_out_1_137;

     reg [1:0] op_in_1_137;
     wire [1:0] op_out_1_137;

     wire r_1_137;

     reg data_in_1_137;
     wire data_out_1_137;

     reg pivot_in_1_137;
     wire pivot_out_1_137;

     always @(posedge clk) begin
         op_in_1_137 <= op_out_1_136;
         pivot_in_1_137 <= pivot_out_1_136;
         start_in_1_137 <= start_out_1_136;
         swap_in_1_137 <= swap_out_1_136;
     end

     always @(posedge clk) begin
         data_in_1_137 <= data_out_0_137;
     end
  
     processor_AB AB_1_137 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_137),
       .start_in   (start_in_1_137),
       .swap_in   (swap_in_1_137),
       .op_in      (op_in_1_137),
       .pivot_in   (pivot_in_1_137),
       .start_out  (start_out_1_137),
       .swap_out   (swap_out_1_137),
       .data_out   (data_out_1_137),
       .op_out     (op_out_1_137),
       .pivot_out  (pivot_out_1_137),
       .r          (r_1_137)
     );

  // row 1, col 138

     reg start_in_1_138;
     wire start_out_1_138;

     reg swap_in_1_138;
     wire swap_out_1_138;

     reg [1:0] op_in_1_138;
     wire [1:0] op_out_1_138;

     wire r_1_138;

     reg data_in_1_138;
     wire data_out_1_138;

     reg pivot_in_1_138;
     wire pivot_out_1_138;

     always @(posedge clk) begin
         op_in_1_138 <= op_out_1_137;
         pivot_in_1_138 <= pivot_out_1_137;
         start_in_1_138 <= start_out_1_137;
         swap_in_1_138 <= swap_out_1_137;
     end

     always @(posedge clk) begin
         data_in_1_138 <= data_out_0_138;
     end
  
     processor_AB AB_1_138 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_138),
       .start_in   (start_in_1_138),
       .swap_in   (swap_in_1_138),
       .op_in      (op_in_1_138),
       .pivot_in   (pivot_in_1_138),
       .start_out  (start_out_1_138),
       .swap_out   (swap_out_1_138),
       .data_out   (data_out_1_138),
       .op_out     (op_out_1_138),
       .pivot_out  (pivot_out_1_138),
       .r          (r_1_138)
     );

  // row 1, col 139

     reg start_in_1_139;
     wire start_out_1_139;

     reg swap_in_1_139;
     wire swap_out_1_139;

     reg [1:0] op_in_1_139;
     wire [1:0] op_out_1_139;

     wire r_1_139;

     reg data_in_1_139;
     wire data_out_1_139;

     reg pivot_in_1_139;
     wire pivot_out_1_139;

     always @(posedge clk) begin
         op_in_1_139 <= op_out_1_138;
         pivot_in_1_139 <= pivot_out_1_138;
         start_in_1_139 <= start_out_1_138;
         swap_in_1_139 <= swap_out_1_138;
     end

     always @(posedge clk) begin
         data_in_1_139 <= data_out_0_139;
     end
  
     processor_AB AB_1_139 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_139),
       .start_in   (start_in_1_139),
       .swap_in   (swap_in_1_139),
       .op_in      (op_in_1_139),
       .pivot_in   (pivot_in_1_139),
       .start_out  (start_out_1_139),
       .swap_out   (swap_out_1_139),
       .data_out   (data_out_1_139),
       .op_out     (op_out_1_139),
       .pivot_out  (pivot_out_1_139),
       .r          (r_1_139)
     );

  // row 1, col 140

     reg start_in_1_140;
     wire start_out_1_140;

     reg swap_in_1_140;
     wire swap_out_1_140;

     reg [1:0] op_in_1_140;
     wire [1:0] op_out_1_140;

     wire r_1_140;

     reg data_in_1_140;
     wire data_out_1_140;

     reg pivot_in_1_140;
     wire pivot_out_1_140;

     always @(posedge clk) begin
         op_in_1_140 <= op_out_1_139;
         pivot_in_1_140 <= pivot_out_1_139;
         start_in_1_140 <= start_out_1_139;
         swap_in_1_140 <= swap_out_1_139;
     end

     always @(posedge clk) begin
         data_in_1_140 <= data_out_0_140;
     end
  
     processor_AB AB_1_140 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_140),
       .start_in   (start_in_1_140),
       .swap_in   (swap_in_1_140),
       .op_in      (op_in_1_140),
       .pivot_in   (pivot_in_1_140),
       .start_out  (start_out_1_140),
       .swap_out   (swap_out_1_140),
       .data_out   (data_out_1_140),
       .op_out     (op_out_1_140),
       .pivot_out  (pivot_out_1_140),
       .r          (r_1_140)
     );

  // row 1, col 141

     reg start_in_1_141;
     wire start_out_1_141;

     reg swap_in_1_141;
     wire swap_out_1_141;

     reg [1:0] op_in_1_141;
     wire [1:0] op_out_1_141;

     wire r_1_141;

     reg data_in_1_141;
     wire data_out_1_141;

     reg pivot_in_1_141;
     wire pivot_out_1_141;

     always @(posedge clk) begin
         op_in_1_141 <= op_out_1_140;
         pivot_in_1_141 <= pivot_out_1_140;
         start_in_1_141 <= start_out_1_140;
         swap_in_1_141 <= swap_out_1_140;
     end

     always @(posedge clk) begin
         data_in_1_141 <= data_out_0_141;
     end
  
     processor_AB AB_1_141 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_141),
       .start_in   (start_in_1_141),
       .swap_in   (swap_in_1_141),
       .op_in      (op_in_1_141),
       .pivot_in   (pivot_in_1_141),
       .start_out  (start_out_1_141),
       .swap_out   (swap_out_1_141),
       .data_out   (data_out_1_141),
       .op_out     (op_out_1_141),
       .pivot_out  (pivot_out_1_141),
       .r          (r_1_141)
     );

  // row 1, col 142

     reg start_in_1_142;
     wire start_out_1_142;

     reg swap_in_1_142;
     wire swap_out_1_142;

     reg [1:0] op_in_1_142;
     wire [1:0] op_out_1_142;

     wire r_1_142;

     reg data_in_1_142;
     wire data_out_1_142;

     reg pivot_in_1_142;
     wire pivot_out_1_142;

     always @(posedge clk) begin
         op_in_1_142 <= op_out_1_141;
         pivot_in_1_142 <= pivot_out_1_141;
         start_in_1_142 <= start_out_1_141;
         swap_in_1_142 <= swap_out_1_141;
     end

     always @(posedge clk) begin
         data_in_1_142 <= data_out_0_142;
     end
  
     processor_AB AB_1_142 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_142),
       .start_in   (start_in_1_142),
       .swap_in   (swap_in_1_142),
       .op_in      (op_in_1_142),
       .pivot_in   (pivot_in_1_142),
       .start_out  (start_out_1_142),
       .swap_out   (swap_out_1_142),
       .data_out   (data_out_1_142),
       .op_out     (op_out_1_142),
       .pivot_out  (pivot_out_1_142),
       .r          (r_1_142)
     );

  // row 1, col 143

     reg start_in_1_143;
     wire start_out_1_143;

     reg swap_in_1_143;
     wire swap_out_1_143;

     reg [1:0] op_in_1_143;
     wire [1:0] op_out_1_143;

     wire r_1_143;

     reg data_in_1_143;
     wire data_out_1_143;

     reg pivot_in_1_143;
     wire pivot_out_1_143;

     always @(posedge clk) begin
         op_in_1_143 <= op_out_1_142;
         pivot_in_1_143 <= pivot_out_1_142;
         start_in_1_143 <= start_out_1_142;
         swap_in_1_143 <= swap_out_1_142;
     end

     always @(posedge clk) begin
         data_in_1_143 <= data_out_0_143;
     end
  
     processor_AB AB_1_143 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_143),
       .start_in   (start_in_1_143),
       .swap_in   (swap_in_1_143),
       .op_in      (op_in_1_143),
       .pivot_in   (pivot_in_1_143),
       .start_out  (start_out_1_143),
       .swap_out   (swap_out_1_143),
       .data_out   (data_out_1_143),
       .op_out     (op_out_1_143),
       .pivot_out  (pivot_out_1_143),
       .r          (r_1_143)
     );

  // row 1, col 144

     reg start_in_1_144;
     wire start_out_1_144;

     reg swap_in_1_144;
     wire swap_out_1_144;

     reg [1:0] op_in_1_144;
     wire [1:0] op_out_1_144;

     wire r_1_144;

     reg data_in_1_144;
     wire data_out_1_144;

     reg pivot_in_1_144;
     wire pivot_out_1_144;

     always @(posedge clk) begin
         op_in_1_144 <= op_out_1_143;
         pivot_in_1_144 <= pivot_out_1_143;
         start_in_1_144 <= start_out_1_143;
         swap_in_1_144 <= swap_out_1_143;
     end

     always @(posedge clk) begin
         data_in_1_144 <= data_out_0_144;
     end
  
     processor_AB AB_1_144 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_144),
       .start_in   (start_in_1_144),
       .swap_in   (swap_in_1_144),
       .op_in      (op_in_1_144),
       .pivot_in   (pivot_in_1_144),
       .start_out  (start_out_1_144),
       .swap_out   (swap_out_1_144),
       .data_out   (data_out_1_144),
       .op_out     (op_out_1_144),
       .pivot_out  (pivot_out_1_144),
       .r          (r_1_144)
     );

  // row 1, col 145

     reg start_in_1_145;
     wire start_out_1_145;

     reg swap_in_1_145;
     wire swap_out_1_145;

     reg [1:0] op_in_1_145;
     wire [1:0] op_out_1_145;

     wire r_1_145;

     reg data_in_1_145;
     wire data_out_1_145;

     reg pivot_in_1_145;
     wire pivot_out_1_145;

     always @(posedge clk) begin
         op_in_1_145 <= op_out_1_144;
         pivot_in_1_145 <= pivot_out_1_144;
         start_in_1_145 <= start_out_1_144;
         swap_in_1_145 <= swap_out_1_144;
     end

     always @(posedge clk) begin
         data_in_1_145 <= data_out_0_145;
     end
  
     processor_AB AB_1_145 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_145),
       .start_in   (start_in_1_145),
       .swap_in   (swap_in_1_145),
       .op_in      (op_in_1_145),
       .pivot_in   (pivot_in_1_145),
       .start_out  (start_out_1_145),
       .swap_out   (swap_out_1_145),
       .data_out   (data_out_1_145),
       .op_out     (op_out_1_145),
       .pivot_out  (pivot_out_1_145),
       .r          (r_1_145)
     );

  // row 1, col 146

     reg start_in_1_146;
     wire start_out_1_146;

     reg swap_in_1_146;
     wire swap_out_1_146;

     reg [1:0] op_in_1_146;
     wire [1:0] op_out_1_146;

     wire r_1_146;

     reg data_in_1_146;
     wire data_out_1_146;

     reg pivot_in_1_146;
     wire pivot_out_1_146;

     always @(posedge clk) begin
         op_in_1_146 <= op_out_1_145;
         pivot_in_1_146 <= pivot_out_1_145;
         start_in_1_146 <= start_out_1_145;
         swap_in_1_146 <= swap_out_1_145;
     end

     always @(posedge clk) begin
         data_in_1_146 <= data_out_0_146;
     end
  
     processor_AB AB_1_146 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_146),
       .start_in   (start_in_1_146),
       .swap_in   (swap_in_1_146),
       .op_in      (op_in_1_146),
       .pivot_in   (pivot_in_1_146),
       .start_out  (start_out_1_146),
       .swap_out   (swap_out_1_146),
       .data_out   (data_out_1_146),
       .op_out     (op_out_1_146),
       .pivot_out  (pivot_out_1_146),
       .r          (r_1_146)
     );

  // row 1, col 147

     reg start_in_1_147;
     wire start_out_1_147;

     reg swap_in_1_147;
     wire swap_out_1_147;

     reg [1:0] op_in_1_147;
     wire [1:0] op_out_1_147;

     wire r_1_147;

     reg data_in_1_147;
     wire data_out_1_147;

     reg pivot_in_1_147;
     wire pivot_out_1_147;

     always @(posedge clk) begin
         op_in_1_147 <= op_out_1_146;
         pivot_in_1_147 <= pivot_out_1_146;
         start_in_1_147 <= start_out_1_146;
         swap_in_1_147 <= swap_out_1_146;
     end

     always @(posedge clk) begin
         data_in_1_147 <= data_out_0_147;
     end
  
     processor_AB AB_1_147 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_147),
       .start_in   (start_in_1_147),
       .swap_in   (swap_in_1_147),
       .op_in      (op_in_1_147),
       .pivot_in   (pivot_in_1_147),
       .start_out  (start_out_1_147),
       .swap_out   (swap_out_1_147),
       .data_out   (data_out_1_147),
       .op_out     (op_out_1_147),
       .pivot_out  (pivot_out_1_147),
       .r          (r_1_147)
     );

  // row 1, col 148

     reg start_in_1_148;
     wire start_out_1_148;

     reg swap_in_1_148;
     wire swap_out_1_148;

     reg [1:0] op_in_1_148;
     wire [1:0] op_out_1_148;

     wire r_1_148;

     reg data_in_1_148;
     wire data_out_1_148;

     reg pivot_in_1_148;
     wire pivot_out_1_148;

     always @(posedge clk) begin
         op_in_1_148 <= op_out_1_147;
         pivot_in_1_148 <= pivot_out_1_147;
         start_in_1_148 <= start_out_1_147;
         swap_in_1_148 <= swap_out_1_147;
     end

     always @(posedge clk) begin
         data_in_1_148 <= data_out_0_148;
     end
  
     processor_AB AB_1_148 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_148),
       .start_in   (start_in_1_148),
       .swap_in   (swap_in_1_148),
       .op_in      (op_in_1_148),
       .pivot_in   (pivot_in_1_148),
       .start_out  (start_out_1_148),
       .swap_out   (swap_out_1_148),
       .data_out   (data_out_1_148),
       .op_out     (op_out_1_148),
       .pivot_out  (pivot_out_1_148),
       .r          (r_1_148)
     );

  // row 1, col 149

     reg start_in_1_149;
     wire start_out_1_149;

     reg swap_in_1_149;
     wire swap_out_1_149;

     reg [1:0] op_in_1_149;
     wire [1:0] op_out_1_149;

     wire r_1_149;

     reg data_in_1_149;
     wire data_out_1_149;

     reg pivot_in_1_149;
     wire pivot_out_1_149;

     always @(posedge clk) begin
         op_in_1_149 <= op_out_1_148;
         pivot_in_1_149 <= pivot_out_1_148;
         start_in_1_149 <= start_out_1_148;
         swap_in_1_149 <= swap_out_1_148;
     end

     always @(posedge clk) begin
         data_in_1_149 <= data_out_0_149;
     end
  
     processor_AB AB_1_149 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_149),
       .start_in   (start_in_1_149),
       .swap_in   (swap_in_1_149),
       .op_in      (op_in_1_149),
       .pivot_in   (pivot_in_1_149),
       .start_out  (start_out_1_149),
       .swap_out   (swap_out_1_149),
       .data_out   (data_out_1_149),
       .op_out     (op_out_1_149),
       .pivot_out  (pivot_out_1_149),
       .r          (r_1_149)
     );

  // row 1, col 150

     reg start_in_1_150;
     wire start_out_1_150;

     reg swap_in_1_150;
     wire swap_out_1_150;

     reg [1:0] op_in_1_150;
     wire [1:0] op_out_1_150;

     wire r_1_150;

     reg data_in_1_150;
     wire data_out_1_150;

     reg pivot_in_1_150;
     wire pivot_out_1_150;

     always @(posedge clk) begin
         op_in_1_150 <= op_out_1_149;
         pivot_in_1_150 <= pivot_out_1_149;
         start_in_1_150 <= start_out_1_149;
         swap_in_1_150 <= swap_out_1_149;
     end

     always @(posedge clk) begin
         data_in_1_150 <= data_out_0_150;
     end
  
     processor_AB AB_1_150 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_150),
       .start_in   (start_in_1_150),
       .swap_in   (swap_in_1_150),
       .op_in      (op_in_1_150),
       .pivot_in   (pivot_in_1_150),
       .start_out  (start_out_1_150),
       .swap_out   (swap_out_1_150),
       .data_out   (data_out_1_150),
       .op_out     (op_out_1_150),
       .pivot_out  (pivot_out_1_150),
       .r          (r_1_150)
     );

  // row 1, col 151

     reg start_in_1_151;
     wire start_out_1_151;

     reg swap_in_1_151;
     wire swap_out_1_151;

     reg [1:0] op_in_1_151;
     wire [1:0] op_out_1_151;

     wire r_1_151;

     reg data_in_1_151;
     wire data_out_1_151;

     reg pivot_in_1_151;
     wire pivot_out_1_151;

     always @(posedge clk) begin
         op_in_1_151 <= op_out_1_150;
         pivot_in_1_151 <= pivot_out_1_150;
         start_in_1_151 <= start_out_1_150;
         swap_in_1_151 <= swap_out_1_150;
     end

     always @(posedge clk) begin
         data_in_1_151 <= data_out_0_151;
     end
  
     processor_AB AB_1_151 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_151),
       .start_in   (start_in_1_151),
       .swap_in   (swap_in_1_151),
       .op_in      (op_in_1_151),
       .pivot_in   (pivot_in_1_151),
       .start_out  (start_out_1_151),
       .swap_out   (swap_out_1_151),
       .data_out   (data_out_1_151),
       .op_out     (op_out_1_151),
       .pivot_out  (pivot_out_1_151),
       .r          (r_1_151)
     );

  // row 1, col 152

     reg start_in_1_152;
     wire start_out_1_152;

     reg swap_in_1_152;
     wire swap_out_1_152;

     reg [1:0] op_in_1_152;
     wire [1:0] op_out_1_152;

     wire r_1_152;

     reg data_in_1_152;
     wire data_out_1_152;

     reg pivot_in_1_152;
     wire pivot_out_1_152;

     always @(posedge clk) begin
         op_in_1_152 <= op_out_1_151;
         pivot_in_1_152 <= pivot_out_1_151;
         start_in_1_152 <= start_out_1_151;
         swap_in_1_152 <= swap_out_1_151;
     end

     always @(posedge clk) begin
         data_in_1_152 <= data_out_0_152;
     end
  
     processor_AB AB_1_152 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_152),
       .start_in   (start_in_1_152),
       .swap_in   (swap_in_1_152),
       .op_in      (op_in_1_152),
       .pivot_in   (pivot_in_1_152),
       .start_out  (start_out_1_152),
       .swap_out   (swap_out_1_152),
       .data_out   (data_out_1_152),
       .op_out     (op_out_1_152),
       .pivot_out  (pivot_out_1_152),
       .r          (r_1_152)
     );

  // row 1, col 153

     reg start_in_1_153;
     wire start_out_1_153;

     reg swap_in_1_153;
     wire swap_out_1_153;

     reg [1:0] op_in_1_153;
     wire [1:0] op_out_1_153;

     wire r_1_153;

     reg data_in_1_153;
     wire data_out_1_153;

     reg pivot_in_1_153;
     wire pivot_out_1_153;

     always @(posedge clk) begin
         op_in_1_153 <= op_out_1_152;
         pivot_in_1_153 <= pivot_out_1_152;
         start_in_1_153 <= start_out_1_152;
         swap_in_1_153 <= swap_out_1_152;
     end

     always @(posedge clk) begin
         data_in_1_153 <= data_out_0_153;
     end
  
     processor_AB AB_1_153 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_153),
       .start_in   (start_in_1_153),
       .swap_in   (swap_in_1_153),
       .op_in      (op_in_1_153),
       .pivot_in   (pivot_in_1_153),
       .start_out  (start_out_1_153),
       .swap_out   (swap_out_1_153),
       .data_out   (data_out_1_153),
       .op_out     (op_out_1_153),
       .pivot_out  (pivot_out_1_153),
       .r          (r_1_153)
     );

  // row 1, col 154

     reg start_in_1_154;
     wire start_out_1_154;

     reg swap_in_1_154;
     wire swap_out_1_154;

     reg [1:0] op_in_1_154;
     wire [1:0] op_out_1_154;

     wire r_1_154;

     reg data_in_1_154;
     wire data_out_1_154;

     reg pivot_in_1_154;
     wire pivot_out_1_154;

     always @(posedge clk) begin
         op_in_1_154 <= op_out_1_153;
         pivot_in_1_154 <= pivot_out_1_153;
         start_in_1_154 <= start_out_1_153;
         swap_in_1_154 <= swap_out_1_153;
     end

     always @(posedge clk) begin
         data_in_1_154 <= data_out_0_154;
     end
  
     processor_AB AB_1_154 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_154),
       .start_in   (start_in_1_154),
       .swap_in   (swap_in_1_154),
       .op_in      (op_in_1_154),
       .pivot_in   (pivot_in_1_154),
       .start_out  (start_out_1_154),
       .swap_out   (swap_out_1_154),
       .data_out   (data_out_1_154),
       .op_out     (op_out_1_154),
       .pivot_out  (pivot_out_1_154),
       .r          (r_1_154)
     );

  // row 1, col 155

     reg start_in_1_155;
     wire start_out_1_155;

     reg swap_in_1_155;
     wire swap_out_1_155;

     reg [1:0] op_in_1_155;
     wire [1:0] op_out_1_155;

     wire r_1_155;

     reg data_in_1_155;
     wire data_out_1_155;

     reg pivot_in_1_155;
     wire pivot_out_1_155;

     always @(posedge clk) begin
         op_in_1_155 <= op_out_1_154;
         pivot_in_1_155 <= pivot_out_1_154;
         start_in_1_155 <= start_out_1_154;
         swap_in_1_155 <= swap_out_1_154;
     end

     always @(posedge clk) begin
         data_in_1_155 <= data_out_0_155;
     end
  
     processor_AB AB_1_155 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_155),
       .start_in   (start_in_1_155),
       .swap_in   (swap_in_1_155),
       .op_in      (op_in_1_155),
       .pivot_in   (pivot_in_1_155),
       .start_out  (start_out_1_155),
       .swap_out   (swap_out_1_155),
       .data_out   (data_out_1_155),
       .op_out     (op_out_1_155),
       .pivot_out  (pivot_out_1_155),
       .r          (r_1_155)
     );

  // row 1, col 156

     reg start_in_1_156;
     wire start_out_1_156;

     reg swap_in_1_156;
     wire swap_out_1_156;

     reg [1:0] op_in_1_156;
     wire [1:0] op_out_1_156;

     wire r_1_156;

     reg data_in_1_156;
     wire data_out_1_156;

     reg pivot_in_1_156;
     wire pivot_out_1_156;

     always @(posedge clk) begin
         op_in_1_156 <= op_out_1_155;
         pivot_in_1_156 <= pivot_out_1_155;
         start_in_1_156 <= start_out_1_155;
         swap_in_1_156 <= swap_out_1_155;
     end

     always @(posedge clk) begin
         data_in_1_156 <= data_out_0_156;
     end
  
     processor_AB AB_1_156 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_156),
       .start_in   (start_in_1_156),
       .swap_in   (swap_in_1_156),
       .op_in      (op_in_1_156),
       .pivot_in   (pivot_in_1_156),
       .start_out  (start_out_1_156),
       .swap_out   (swap_out_1_156),
       .data_out   (data_out_1_156),
       .op_out     (op_out_1_156),
       .pivot_out  (pivot_out_1_156),
       .r          (r_1_156)
     );

  // row 1, col 157

     reg start_in_1_157;
     wire start_out_1_157;

     reg swap_in_1_157;
     wire swap_out_1_157;

     reg [1:0] op_in_1_157;
     wire [1:0] op_out_1_157;

     wire r_1_157;

     reg data_in_1_157;
     wire data_out_1_157;

     reg pivot_in_1_157;
     wire pivot_out_1_157;

     always @(posedge clk) begin
         op_in_1_157 <= op_out_1_156;
         pivot_in_1_157 <= pivot_out_1_156;
         start_in_1_157 <= start_out_1_156;
         swap_in_1_157 <= swap_out_1_156;
     end

     always @(posedge clk) begin
         data_in_1_157 <= data_out_0_157;
     end
  
     processor_AB AB_1_157 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_157),
       .start_in   (start_in_1_157),
       .swap_in   (swap_in_1_157),
       .op_in      (op_in_1_157),
       .pivot_in   (pivot_in_1_157),
       .start_out  (start_out_1_157),
       .swap_out   (swap_out_1_157),
       .data_out   (data_out_1_157),
       .op_out     (op_out_1_157),
       .pivot_out  (pivot_out_1_157),
       .r          (r_1_157)
     );

  // row 1, col 158

     reg start_in_1_158;
     wire start_out_1_158;

     reg swap_in_1_158;
     wire swap_out_1_158;

     reg [1:0] op_in_1_158;
     wire [1:0] op_out_1_158;

     wire r_1_158;

     reg data_in_1_158;
     wire data_out_1_158;

     reg pivot_in_1_158;
     wire pivot_out_1_158;

     always @(posedge clk) begin
         op_in_1_158 <= op_out_1_157;
         pivot_in_1_158 <= pivot_out_1_157;
         start_in_1_158 <= start_out_1_157;
         swap_in_1_158 <= swap_out_1_157;
     end

     always @(posedge clk) begin
         data_in_1_158 <= data_out_0_158;
     end
  
     processor_AB AB_1_158 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_158),
       .start_in   (start_in_1_158),
       .swap_in   (swap_in_1_158),
       .op_in      (op_in_1_158),
       .pivot_in   (pivot_in_1_158),
       .start_out  (start_out_1_158),
       .swap_out   (swap_out_1_158),
       .data_out   (data_out_1_158),
       .op_out     (op_out_1_158),
       .pivot_out  (pivot_out_1_158),
       .r          (r_1_158)
     );

  // row 1, col 159

     reg start_in_1_159;
     wire start_out_1_159;

     reg swap_in_1_159;
     wire swap_out_1_159;

     reg [1:0] op_in_1_159;
     wire [1:0] op_out_1_159;

     wire r_1_159;

     reg data_in_1_159;
     wire data_out_1_159;

     reg pivot_in_1_159;
     wire pivot_out_1_159;

     always @(posedge clk) begin
         op_in_1_159 <= op_out_1_158;
         pivot_in_1_159 <= pivot_out_1_158;
         start_in_1_159 <= start_out_1_158;
         swap_in_1_159 <= swap_out_1_158;
     end

     always @(posedge clk) begin
         data_in_1_159 <= data_out_0_159;
     end
  
     processor_AB AB_1_159 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_159),
       .start_in   (start_in_1_159),
       .swap_in   (swap_in_1_159),
       .op_in      (op_in_1_159),
       .pivot_in   (pivot_in_1_159),
       .start_out  (start_out_1_159),
       .swap_out   (swap_out_1_159),
       .data_out   (data_out_1_159),
       .op_out     (op_out_1_159),
       .pivot_out  (pivot_out_1_159),
       .r          (r_1_159)
     );

  // row 1, col 160

     reg start_in_1_160;
     wire start_out_1_160;

     reg swap_in_1_160;
     wire swap_out_1_160;

     reg [1:0] op_in_1_160;
     wire [1:0] op_out_1_160;

     wire r_1_160;

     reg data_in_1_160;
     wire data_out_1_160;

     reg pivot_in_1_160;
     wire pivot_out_1_160;

     always @(posedge clk) begin
         op_in_1_160 <= op_out_1_159;
         pivot_in_1_160 <= pivot_out_1_159;
         start_in_1_160 <= start_out_1_159;
         swap_in_1_160 <= swap_out_1_159;
     end

     always @(posedge clk) begin
         data_in_1_160 <= data_out_0_160;
     end
  
     processor_AB AB_1_160 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_160),
       .start_in   (start_in_1_160),
       .swap_in   (swap_in_1_160),
       .op_in      (op_in_1_160),
       .pivot_in   (pivot_in_1_160),
       .start_out  (start_out_1_160),
       .swap_out   (swap_out_1_160),
       .data_out   (data_out_1_160),
       .op_out     (op_out_1_160),
       .pivot_out  (pivot_out_1_160),
       .r          (r_1_160)
     );

  // row 1, col 161

     reg start_in_1_161;
     wire start_out_1_161;

     reg swap_in_1_161;
     wire swap_out_1_161;

     reg [1:0] op_in_1_161;
     wire [1:0] op_out_1_161;

     wire r_1_161;

     reg data_in_1_161;
     wire data_out_1_161;

     reg pivot_in_1_161;
     wire pivot_out_1_161;

     always @(posedge clk) begin
         op_in_1_161 <= op_out_1_160;
         pivot_in_1_161 <= pivot_out_1_160;
         start_in_1_161 <= start_out_1_160;
         swap_in_1_161 <= swap_out_1_160;
     end

     always @(posedge clk) begin
         data_in_1_161 <= data_out_0_161;
     end
  
     processor_AB AB_1_161 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_161),
       .start_in   (start_in_1_161),
       .swap_in   (swap_in_1_161),
       .op_in      (op_in_1_161),
       .pivot_in   (pivot_in_1_161),
       .start_out  (start_out_1_161),
       .swap_out   (swap_out_1_161),
       .data_out   (data_out_1_161),
       .op_out     (op_out_1_161),
       .pivot_out  (pivot_out_1_161),
       .r          (r_1_161)
     );

  // row 1, col 162

     reg start_in_1_162;
     wire start_out_1_162;

     reg swap_in_1_162;
     wire swap_out_1_162;

     reg [1:0] op_in_1_162;
     wire [1:0] op_out_1_162;

     wire r_1_162;

     reg data_in_1_162;
     wire data_out_1_162;

     reg pivot_in_1_162;
     wire pivot_out_1_162;

     always @(posedge clk) begin
         op_in_1_162 <= op_out_1_161;
         pivot_in_1_162 <= pivot_out_1_161;
         start_in_1_162 <= start_out_1_161;
         swap_in_1_162 <= swap_out_1_161;
     end

     always @(posedge clk) begin
         data_in_1_162 <= data_out_0_162;
     end
  
     processor_AB AB_1_162 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_162),
       .start_in   (start_in_1_162),
       .swap_in   (swap_in_1_162),
       .op_in      (op_in_1_162),
       .pivot_in   (pivot_in_1_162),
       .start_out  (start_out_1_162),
       .swap_out   (swap_out_1_162),
       .data_out   (data_out_1_162),
       .op_out     (op_out_1_162),
       .pivot_out  (pivot_out_1_162),
       .r          (r_1_162)
     );

  // row 1, col 163

     reg start_in_1_163;
     wire start_out_1_163;

     reg swap_in_1_163;
     wire swap_out_1_163;

     reg [1:0] op_in_1_163;
     wire [1:0] op_out_1_163;

     wire r_1_163;

     reg data_in_1_163;
     wire data_out_1_163;

     reg pivot_in_1_163;
     wire pivot_out_1_163;

     always @(posedge clk) begin
         op_in_1_163 <= op_out_1_162;
         pivot_in_1_163 <= pivot_out_1_162;
         start_in_1_163 <= start_out_1_162;
         swap_in_1_163 <= swap_out_1_162;
     end

     always @(posedge clk) begin
         data_in_1_163 <= data_out_0_163;
     end
  
     processor_AB AB_1_163 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_163),
       .start_in   (start_in_1_163),
       .swap_in   (swap_in_1_163),
       .op_in      (op_in_1_163),
       .pivot_in   (pivot_in_1_163),
       .start_out  (start_out_1_163),
       .swap_out   (swap_out_1_163),
       .data_out   (data_out_1_163),
       .op_out     (op_out_1_163),
       .pivot_out  (pivot_out_1_163),
       .r          (r_1_163)
     );

  // row 1, col 164

     reg start_in_1_164;
     wire start_out_1_164;

     reg swap_in_1_164;
     wire swap_out_1_164;

     reg [1:0] op_in_1_164;
     wire [1:0] op_out_1_164;

     wire r_1_164;

     reg data_in_1_164;
     wire data_out_1_164;

     reg pivot_in_1_164;
     wire pivot_out_1_164;

     always @(posedge clk) begin
         op_in_1_164 <= op_out_1_163;
         pivot_in_1_164 <= pivot_out_1_163;
         start_in_1_164 <= start_out_1_163;
         swap_in_1_164 <= swap_out_1_163;
     end

     always @(posedge clk) begin
         data_in_1_164 <= data_out_0_164;
     end
  
     processor_AB AB_1_164 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_164),
       .start_in   (start_in_1_164),
       .swap_in   (swap_in_1_164),
       .op_in      (op_in_1_164),
       .pivot_in   (pivot_in_1_164),
       .start_out  (start_out_1_164),
       .swap_out   (swap_out_1_164),
       .data_out   (data_out_1_164),
       .op_out     (op_out_1_164),
       .pivot_out  (pivot_out_1_164),
       .r          (r_1_164)
     );

  // row 1, col 165

     reg start_in_1_165;
     wire start_out_1_165;

     reg swap_in_1_165;
     wire swap_out_1_165;

     reg [1:0] op_in_1_165;
     wire [1:0] op_out_1_165;

     wire r_1_165;

     reg data_in_1_165;
     wire data_out_1_165;

     reg pivot_in_1_165;
     wire pivot_out_1_165;

     always @(posedge clk) begin
         op_in_1_165 <= op_out_1_164;
         pivot_in_1_165 <= pivot_out_1_164;
         start_in_1_165 <= start_out_1_164;
         swap_in_1_165 <= swap_out_1_164;
     end

     always @(posedge clk) begin
         data_in_1_165 <= data_out_0_165;
     end
  
     processor_AB AB_1_165 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_1_165),
       .start_in   (start_in_1_165),
       .swap_in   (swap_in_1_165),
       .op_in      (op_in_1_165),
       .pivot_in   (pivot_in_1_165),
       .start_out  (start_out_1_165),
       .swap_out   (swap_out_1_165),
       .data_out   (data_out_1_165),
       .op_out     (op_out_1_165),
       .pivot_out  (pivot_out_1_165),
       .r          (r_1_165)
     );

  /////////////////////////////////////
  // row 2
  // row 2, col 0

     wire start_in_2_0;
     wire start_out_2_0;

     wire swap_in_2_0;
     wire swap_out_2_0;

     wire [1:0] op_in_2_0;
     wire [1:0] op_out_2_0;

     wire r_2_0;

     reg data_in_2_0;
     wire data_out_2_0;

     wire pivot_in_2_0;
     wire pivout_out_2_0;

     assign op_in_2_0 = 2'b00;
     assign pivot_in_2_0 = 0;

     assign start_in_2_0 = start_row[2]; 
     assign swap_in_2_0 = mode ? swap : swap_row[2]; 

     always @(posedge clk) begin
         data_in_2_0 <= data_out_1_0;
     end

     processor_AB AB_2_0 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_0),
       .start_in   (start_in_2_0),
       .swap_in   (swap_in_2_0),
       .op_in      (op_in_2_0),
       .pivot_in   (pivot_in_2_0),
       .start_out  (start_out_2_0),
       .swap_out   (swap_out_2_0),
       .data_out   (data_out_2_0),
       .op_out     (op_out_2_0),
       .pivot_out  (pivot_out_2_0),
       .r          (r_2_0)
     );

  // row 2, col 1

     reg start_in_2_1;
     wire start_out_2_1;

     reg swap_in_2_1;
     wire swap_out_2_1;

     reg [1:0] op_in_2_1;
     wire [1:0] op_out_2_1;

     wire r_2_1;

     reg data_in_2_1;
     wire data_out_2_1;

     reg pivot_in_2_1;
     wire pivot_out_2_1;

     always @(posedge clk) begin
         op_in_2_1 <= op_out_2_0;
         pivot_in_2_1 <= pivot_out_2_0;
         start_in_2_1 <= start_out_2_0;
         swap_in_2_1 <= swap_out_2_0;
     end

     always @(posedge clk) begin
         data_in_2_1 <= data_out_1_1;
     end
  
     processor_AB AB_2_1 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_1),
       .start_in   (start_in_2_1),
       .swap_in   (swap_in_2_1),
       .op_in      (op_in_2_1),
       .pivot_in   (pivot_in_2_1),
       .start_out  (start_out_2_1),
       .swap_out   (swap_out_2_1),
       .data_out   (data_out_2_1),
       .op_out     (op_out_2_1),
       .pivot_out  (pivot_out_2_1),
       .r          (r_2_1)
     );

  // row 2, col 2

     reg start_in_2_2;
     wire start_out_2_2;

     reg swap_in_2_2;
     wire swap_out_2_2;

     reg [1:0] op_in_2_2;
     wire [1:0] op_out_2_2;

     wire r_2_2;

     reg data_in_2_2;
     wire data_out_2_2;

     reg pivot_in_2_2;
     wire pivot_out_2_2;

     always @(posedge clk) begin
         op_in_2_2 <= op_out_2_1;
         pivot_in_2_2 <= pivot_out_2_1;
         start_in_2_2 <= start_out_2_1;
         swap_in_2_2 <= swap_out_2_1;
     end

     always @(posedge clk) begin
         data_in_2_2 <= data_out_1_2;
     end
  
     processor_AB AB_2_2 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_2),
       .start_in   (start_in_2_2),
       .swap_in   (swap_in_2_2),
       .op_in      (op_in_2_2),
       .pivot_in   (pivot_in_2_2),
       .start_out  (start_out_2_2),
       .swap_out   (swap_out_2_2),
       .data_out   (data_out_2_2),
       .op_out     (op_out_2_2),
       .pivot_out  (pivot_out_2_2),
       .r          (r_2_2)
     );

  // row 2, col 3

     reg start_in_2_3;
     wire start_out_2_3;

     reg swap_in_2_3;
     wire swap_out_2_3;

     reg [1:0] op_in_2_3;
     wire [1:0] op_out_2_3;

     wire r_2_3;

     reg data_in_2_3;
     wire data_out_2_3;

     reg pivot_in_2_3;
     wire pivot_out_2_3;

     always @(posedge clk) begin
         op_in_2_3 <= op_out_2_2;
         pivot_in_2_3 <= pivot_out_2_2;
         start_in_2_3 <= start_out_2_2;
         swap_in_2_3 <= swap_out_2_2;
     end

     always @(posedge clk) begin
         data_in_2_3 <= data_out_1_3;
     end
  
     processor_AB AB_2_3 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_3),
       .start_in   (start_in_2_3),
       .swap_in   (swap_in_2_3),
       .op_in      (op_in_2_3),
       .pivot_in   (pivot_in_2_3),
       .start_out  (start_out_2_3),
       .swap_out   (swap_out_2_3),
       .data_out   (data_out_2_3),
       .op_out     (op_out_2_3),
       .pivot_out  (pivot_out_2_3),
       .r          (r_2_3)
     );

  // row 2, col 4

     reg start_in_2_4;
     wire start_out_2_4;

     reg swap_in_2_4;
     wire swap_out_2_4;

     reg [1:0] op_in_2_4;
     wire [1:0] op_out_2_4;

     wire r_2_4;

     reg data_in_2_4;
     wire data_out_2_4;

     reg pivot_in_2_4;
     wire pivot_out_2_4;

     always @(posedge clk) begin
         op_in_2_4 <= op_out_2_3;
         pivot_in_2_4 <= pivot_out_2_3;
         start_in_2_4 <= start_out_2_3;
         swap_in_2_4 <= swap_out_2_3;
     end

     always @(posedge clk) begin
         data_in_2_4 <= data_out_1_4;
     end
  
     processor_AB AB_2_4 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_4),
       .start_in   (start_in_2_4),
       .swap_in   (swap_in_2_4),
       .op_in      (op_in_2_4),
       .pivot_in   (pivot_in_2_4),
       .start_out  (start_out_2_4),
       .swap_out   (swap_out_2_4),
       .data_out   (data_out_2_4),
       .op_out     (op_out_2_4),
       .pivot_out  (pivot_out_2_4),
       .r          (r_2_4)
     );

  // row 2, col 5

     reg start_in_2_5;
     wire start_out_2_5;

     reg swap_in_2_5;
     wire swap_out_2_5;

     reg [1:0] op_in_2_5;
     wire [1:0] op_out_2_5;

     wire r_2_5;

     reg data_in_2_5;
     wire data_out_2_5;

     reg pivot_in_2_5;
     wire pivot_out_2_5;

     always @(posedge clk) begin
         op_in_2_5 <= op_out_2_4;
         pivot_in_2_5 <= pivot_out_2_4;
         start_in_2_5 <= start_out_2_4;
         swap_in_2_5 <= swap_out_2_4;
     end

     always @(posedge clk) begin
         data_in_2_5 <= data_out_1_5;
     end
  
     processor_AB AB_2_5 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_5),
       .start_in   (start_in_2_5),
       .swap_in   (swap_in_2_5),
       .op_in      (op_in_2_5),
       .pivot_in   (pivot_in_2_5),
       .start_out  (start_out_2_5),
       .swap_out   (swap_out_2_5),
       .data_out   (data_out_2_5),
       .op_out     (op_out_2_5),
       .pivot_out  (pivot_out_2_5),
       .r          (r_2_5)
     );

  // row 2, col 6

     reg start_in_2_6;
     wire start_out_2_6;

     reg swap_in_2_6;
     wire swap_out_2_6;

     reg [1:0] op_in_2_6;
     wire [1:0] op_out_2_6;

     wire r_2_6;

     reg data_in_2_6;
     wire data_out_2_6;

     reg pivot_in_2_6;
     wire pivot_out_2_6;

     always @(posedge clk) begin
         op_in_2_6 <= op_out_2_5;
         pivot_in_2_6 <= pivot_out_2_5;
         start_in_2_6 <= start_out_2_5;
         swap_in_2_6 <= swap_out_2_5;
     end

     always @(posedge clk) begin
         data_in_2_6 <= data_out_1_6;
     end
  
     processor_AB AB_2_6 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_6),
       .start_in   (start_in_2_6),
       .swap_in   (swap_in_2_6),
       .op_in      (op_in_2_6),
       .pivot_in   (pivot_in_2_6),
       .start_out  (start_out_2_6),
       .swap_out   (swap_out_2_6),
       .data_out   (data_out_2_6),
       .op_out     (op_out_2_6),
       .pivot_out  (pivot_out_2_6),
       .r          (r_2_6)
     );

  // row 2, col 7

     reg start_in_2_7;
     wire start_out_2_7;

     reg swap_in_2_7;
     wire swap_out_2_7;

     reg [1:0] op_in_2_7;
     wire [1:0] op_out_2_7;

     wire r_2_7;

     reg data_in_2_7;
     wire data_out_2_7;

     reg pivot_in_2_7;
     wire pivot_out_2_7;

     always @(posedge clk) begin
         op_in_2_7 <= op_out_2_6;
         pivot_in_2_7 <= pivot_out_2_6;
         start_in_2_7 <= start_out_2_6;
         swap_in_2_7 <= swap_out_2_6;
     end

     always @(posedge clk) begin
         data_in_2_7 <= data_out_1_7;
     end
  
     processor_AB AB_2_7 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_7),
       .start_in   (start_in_2_7),
       .swap_in   (swap_in_2_7),
       .op_in      (op_in_2_7),
       .pivot_in   (pivot_in_2_7),
       .start_out  (start_out_2_7),
       .swap_out   (swap_out_2_7),
       .data_out   (data_out_2_7),
       .op_out     (op_out_2_7),
       .pivot_out  (pivot_out_2_7),
       .r          (r_2_7)
     );

  // row 2, col 8

     reg start_in_2_8;
     wire start_out_2_8;

     reg swap_in_2_8;
     wire swap_out_2_8;

     reg [1:0] op_in_2_8;
     wire [1:0] op_out_2_8;

     wire r_2_8;

     reg data_in_2_8;
     wire data_out_2_8;

     reg pivot_in_2_8;
     wire pivot_out_2_8;

     always @(posedge clk) begin
         op_in_2_8 <= op_out_2_7;
         pivot_in_2_8 <= pivot_out_2_7;
         start_in_2_8 <= start_out_2_7;
         swap_in_2_8 <= swap_out_2_7;
     end

     always @(posedge clk) begin
         data_in_2_8 <= data_out_1_8;
     end
  
     processor_AB AB_2_8 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_8),
       .start_in   (start_in_2_8),
       .swap_in   (swap_in_2_8),
       .op_in      (op_in_2_8),
       .pivot_in   (pivot_in_2_8),
       .start_out  (start_out_2_8),
       .swap_out   (swap_out_2_8),
       .data_out   (data_out_2_8),
       .op_out     (op_out_2_8),
       .pivot_out  (pivot_out_2_8),
       .r          (r_2_8)
     );

  // row 2, col 9

     reg start_in_2_9;
     wire start_out_2_9;

     reg swap_in_2_9;
     wire swap_out_2_9;

     reg [1:0] op_in_2_9;
     wire [1:0] op_out_2_9;

     wire r_2_9;

     reg data_in_2_9;
     wire data_out_2_9;

     reg pivot_in_2_9;
     wire pivot_out_2_9;

     always @(posedge clk) begin
         op_in_2_9 <= op_out_2_8;
         pivot_in_2_9 <= pivot_out_2_8;
         start_in_2_9 <= start_out_2_8;
         swap_in_2_9 <= swap_out_2_8;
     end

     always @(posedge clk) begin
         data_in_2_9 <= data_out_1_9;
     end
  
     processor_AB AB_2_9 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_9),
       .start_in   (start_in_2_9),
       .swap_in   (swap_in_2_9),
       .op_in      (op_in_2_9),
       .pivot_in   (pivot_in_2_9),
       .start_out  (start_out_2_9),
       .swap_out   (swap_out_2_9),
       .data_out   (data_out_2_9),
       .op_out     (op_out_2_9),
       .pivot_out  (pivot_out_2_9),
       .r          (r_2_9)
     );

  // row 2, col 10

     reg start_in_2_10;
     wire start_out_2_10;

     reg swap_in_2_10;
     wire swap_out_2_10;

     reg [1:0] op_in_2_10;
     wire [1:0] op_out_2_10;

     wire r_2_10;

     reg data_in_2_10;
     wire data_out_2_10;

     reg pivot_in_2_10;
     wire pivot_out_2_10;

     always @(posedge clk) begin
         op_in_2_10 <= op_out_2_9;
         pivot_in_2_10 <= pivot_out_2_9;
         start_in_2_10 <= start_out_2_9;
         swap_in_2_10 <= swap_out_2_9;
     end

     always @(posedge clk) begin
         data_in_2_10 <= data_out_1_10;
     end
  
     processor_AB AB_2_10 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_10),
       .start_in   (start_in_2_10),
       .swap_in   (swap_in_2_10),
       .op_in      (op_in_2_10),
       .pivot_in   (pivot_in_2_10),
       .start_out  (start_out_2_10),
       .swap_out   (swap_out_2_10),
       .data_out   (data_out_2_10),
       .op_out     (op_out_2_10),
       .pivot_out  (pivot_out_2_10),
       .r          (r_2_10)
     );

  // row 2, col 11

     reg start_in_2_11;
     wire start_out_2_11;

     reg swap_in_2_11;
     wire swap_out_2_11;

     reg [1:0] op_in_2_11;
     wire [1:0] op_out_2_11;

     wire r_2_11;

     reg data_in_2_11;
     wire data_out_2_11;

     reg pivot_in_2_11;
     wire pivot_out_2_11;

     always @(posedge clk) begin
         op_in_2_11 <= op_out_2_10;
         pivot_in_2_11 <= pivot_out_2_10;
         start_in_2_11 <= start_out_2_10;
         swap_in_2_11 <= swap_out_2_10;
     end

     always @(posedge clk) begin
         data_in_2_11 <= data_out_1_11;
     end
  
     processor_AB AB_2_11 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_11),
       .start_in   (start_in_2_11),
       .swap_in   (swap_in_2_11),
       .op_in      (op_in_2_11),
       .pivot_in   (pivot_in_2_11),
       .start_out  (start_out_2_11),
       .swap_out   (swap_out_2_11),
       .data_out   (data_out_2_11),
       .op_out     (op_out_2_11),
       .pivot_out  (pivot_out_2_11),
       .r          (r_2_11)
     );

  // row 2, col 12

     reg start_in_2_12;
     wire start_out_2_12;

     reg swap_in_2_12;
     wire swap_out_2_12;

     reg [1:0] op_in_2_12;
     wire [1:0] op_out_2_12;

     wire r_2_12;

     reg data_in_2_12;
     wire data_out_2_12;

     reg pivot_in_2_12;
     wire pivot_out_2_12;

     always @(posedge clk) begin
         op_in_2_12 <= op_out_2_11;
         pivot_in_2_12 <= pivot_out_2_11;
         start_in_2_12 <= start_out_2_11;
         swap_in_2_12 <= swap_out_2_11;
     end

     always @(posedge clk) begin
         data_in_2_12 <= data_out_1_12;
     end
  
     processor_AB AB_2_12 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_12),
       .start_in   (start_in_2_12),
       .swap_in   (swap_in_2_12),
       .op_in      (op_in_2_12),
       .pivot_in   (pivot_in_2_12),
       .start_out  (start_out_2_12),
       .swap_out   (swap_out_2_12),
       .data_out   (data_out_2_12),
       .op_out     (op_out_2_12),
       .pivot_out  (pivot_out_2_12),
       .r          (r_2_12)
     );

  // row 2, col 13

     reg start_in_2_13;
     wire start_out_2_13;

     reg swap_in_2_13;
     wire swap_out_2_13;

     reg [1:0] op_in_2_13;
     wire [1:0] op_out_2_13;

     wire r_2_13;

     reg data_in_2_13;
     wire data_out_2_13;

     reg pivot_in_2_13;
     wire pivot_out_2_13;

     always @(posedge clk) begin
         op_in_2_13 <= op_out_2_12;
         pivot_in_2_13 <= pivot_out_2_12;
         start_in_2_13 <= start_out_2_12;
         swap_in_2_13 <= swap_out_2_12;
     end

     always @(posedge clk) begin
         data_in_2_13 <= data_out_1_13;
     end
  
     processor_AB AB_2_13 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_13),
       .start_in   (start_in_2_13),
       .swap_in   (swap_in_2_13),
       .op_in      (op_in_2_13),
       .pivot_in   (pivot_in_2_13),
       .start_out  (start_out_2_13),
       .swap_out   (swap_out_2_13),
       .data_out   (data_out_2_13),
       .op_out     (op_out_2_13),
       .pivot_out  (pivot_out_2_13),
       .r          (r_2_13)
     );

  // row 2, col 14

     reg start_in_2_14;
     wire start_out_2_14;

     reg swap_in_2_14;
     wire swap_out_2_14;

     reg [1:0] op_in_2_14;
     wire [1:0] op_out_2_14;

     wire r_2_14;

     reg data_in_2_14;
     wire data_out_2_14;

     reg pivot_in_2_14;
     wire pivot_out_2_14;

     always @(posedge clk) begin
         op_in_2_14 <= op_out_2_13;
         pivot_in_2_14 <= pivot_out_2_13;
         start_in_2_14 <= start_out_2_13;
         swap_in_2_14 <= swap_out_2_13;
     end

     always @(posedge clk) begin
         data_in_2_14 <= data_out_1_14;
     end
  
     processor_AB AB_2_14 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_14),
       .start_in   (start_in_2_14),
       .swap_in   (swap_in_2_14),
       .op_in      (op_in_2_14),
       .pivot_in   (pivot_in_2_14),
       .start_out  (start_out_2_14),
       .swap_out   (swap_out_2_14),
       .data_out   (data_out_2_14),
       .op_out     (op_out_2_14),
       .pivot_out  (pivot_out_2_14),
       .r          (r_2_14)
     );

  // row 2, col 15

     reg start_in_2_15;
     wire start_out_2_15;

     reg swap_in_2_15;
     wire swap_out_2_15;

     reg [1:0] op_in_2_15;
     wire [1:0] op_out_2_15;

     wire r_2_15;

     reg data_in_2_15;
     wire data_out_2_15;

     reg pivot_in_2_15;
     wire pivot_out_2_15;

     always @(posedge clk) begin
         op_in_2_15 <= op_out_2_14;
         pivot_in_2_15 <= pivot_out_2_14;
         start_in_2_15 <= start_out_2_14;
         swap_in_2_15 <= swap_out_2_14;
     end

     always @(posedge clk) begin
         data_in_2_15 <= data_out_1_15;
     end
  
     processor_AB AB_2_15 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_15),
       .start_in   (start_in_2_15),
       .swap_in   (swap_in_2_15),
       .op_in      (op_in_2_15),
       .pivot_in   (pivot_in_2_15),
       .start_out  (start_out_2_15),
       .swap_out   (swap_out_2_15),
       .data_out   (data_out_2_15),
       .op_out     (op_out_2_15),
       .pivot_out  (pivot_out_2_15),
       .r          (r_2_15)
     );

  // row 2, col 16

     reg start_in_2_16;
     wire start_out_2_16;

     reg swap_in_2_16;
     wire swap_out_2_16;

     reg [1:0] op_in_2_16;
     wire [1:0] op_out_2_16;

     wire r_2_16;

     reg data_in_2_16;
     wire data_out_2_16;

     reg pivot_in_2_16;
     wire pivot_out_2_16;

     always @(posedge clk) begin
         op_in_2_16 <= op_out_2_15;
         pivot_in_2_16 <= pivot_out_2_15;
         start_in_2_16 <= start_out_2_15;
         swap_in_2_16 <= swap_out_2_15;
     end

     always @(posedge clk) begin
         data_in_2_16 <= data_out_1_16;
     end
  
     processor_AB AB_2_16 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_16),
       .start_in   (start_in_2_16),
       .swap_in   (swap_in_2_16),
       .op_in      (op_in_2_16),
       .pivot_in   (pivot_in_2_16),
       .start_out  (start_out_2_16),
       .swap_out   (swap_out_2_16),
       .data_out   (data_out_2_16),
       .op_out     (op_out_2_16),
       .pivot_out  (pivot_out_2_16),
       .r          (r_2_16)
     );

  // row 2, col 17

     reg start_in_2_17;
     wire start_out_2_17;

     reg swap_in_2_17;
     wire swap_out_2_17;

     reg [1:0] op_in_2_17;
     wire [1:0] op_out_2_17;

     wire r_2_17;

     reg data_in_2_17;
     wire data_out_2_17;

     reg pivot_in_2_17;
     wire pivot_out_2_17;

     always @(posedge clk) begin
         op_in_2_17 <= op_out_2_16;
         pivot_in_2_17 <= pivot_out_2_16;
         start_in_2_17 <= start_out_2_16;
         swap_in_2_17 <= swap_out_2_16;
     end

     always @(posedge clk) begin
         data_in_2_17 <= data_out_1_17;
     end
  
     processor_AB AB_2_17 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_17),
       .start_in   (start_in_2_17),
       .swap_in   (swap_in_2_17),
       .op_in      (op_in_2_17),
       .pivot_in   (pivot_in_2_17),
       .start_out  (start_out_2_17),
       .swap_out   (swap_out_2_17),
       .data_out   (data_out_2_17),
       .op_out     (op_out_2_17),
       .pivot_out  (pivot_out_2_17),
       .r          (r_2_17)
     );

  // row 2, col 18

     reg start_in_2_18;
     wire start_out_2_18;

     reg swap_in_2_18;
     wire swap_out_2_18;

     reg [1:0] op_in_2_18;
     wire [1:0] op_out_2_18;

     wire r_2_18;

     reg data_in_2_18;
     wire data_out_2_18;

     reg pivot_in_2_18;
     wire pivot_out_2_18;

     always @(posedge clk) begin
         op_in_2_18 <= op_out_2_17;
         pivot_in_2_18 <= pivot_out_2_17;
         start_in_2_18 <= start_out_2_17;
         swap_in_2_18 <= swap_out_2_17;
     end

     always @(posedge clk) begin
         data_in_2_18 <= data_out_1_18;
     end
  
     processor_AB AB_2_18 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_18),
       .start_in   (start_in_2_18),
       .swap_in   (swap_in_2_18),
       .op_in      (op_in_2_18),
       .pivot_in   (pivot_in_2_18),
       .start_out  (start_out_2_18),
       .swap_out   (swap_out_2_18),
       .data_out   (data_out_2_18),
       .op_out     (op_out_2_18),
       .pivot_out  (pivot_out_2_18),
       .r          (r_2_18)
     );

  // row 2, col 19

     reg start_in_2_19;
     wire start_out_2_19;

     reg swap_in_2_19;
     wire swap_out_2_19;

     reg [1:0] op_in_2_19;
     wire [1:0] op_out_2_19;

     wire r_2_19;

     reg data_in_2_19;
     wire data_out_2_19;

     reg pivot_in_2_19;
     wire pivot_out_2_19;

     always @(posedge clk) begin
         op_in_2_19 <= op_out_2_18;
         pivot_in_2_19 <= pivot_out_2_18;
         start_in_2_19 <= start_out_2_18;
         swap_in_2_19 <= swap_out_2_18;
     end

     always @(posedge clk) begin
         data_in_2_19 <= data_out_1_19;
     end
  
     processor_AB AB_2_19 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_19),
       .start_in   (start_in_2_19),
       .swap_in   (swap_in_2_19),
       .op_in      (op_in_2_19),
       .pivot_in   (pivot_in_2_19),
       .start_out  (start_out_2_19),
       .swap_out   (swap_out_2_19),
       .data_out   (data_out_2_19),
       .op_out     (op_out_2_19),
       .pivot_out  (pivot_out_2_19),
       .r          (r_2_19)
     );

  // row 2, col 20

     reg start_in_2_20;
     wire start_out_2_20;

     reg swap_in_2_20;
     wire swap_out_2_20;

     reg [1:0] op_in_2_20;
     wire [1:0] op_out_2_20;

     wire r_2_20;

     reg data_in_2_20;
     wire data_out_2_20;

     reg pivot_in_2_20;
     wire pivot_out_2_20;

     always @(posedge clk) begin
         op_in_2_20 <= op_out_2_19;
         pivot_in_2_20 <= pivot_out_2_19;
         start_in_2_20 <= start_out_2_19;
         swap_in_2_20 <= swap_out_2_19;
     end

     always @(posedge clk) begin
         data_in_2_20 <= data_out_1_20;
     end
  
     processor_AB AB_2_20 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_20),
       .start_in   (start_in_2_20),
       .swap_in   (swap_in_2_20),
       .op_in      (op_in_2_20),
       .pivot_in   (pivot_in_2_20),
       .start_out  (start_out_2_20),
       .swap_out   (swap_out_2_20),
       .data_out   (data_out_2_20),
       .op_out     (op_out_2_20),
       .pivot_out  (pivot_out_2_20),
       .r          (r_2_20)
     );

  // row 2, col 21

     reg start_in_2_21;
     wire start_out_2_21;

     reg swap_in_2_21;
     wire swap_out_2_21;

     reg [1:0] op_in_2_21;
     wire [1:0] op_out_2_21;

     wire r_2_21;

     reg data_in_2_21;
     wire data_out_2_21;

     reg pivot_in_2_21;
     wire pivot_out_2_21;

     always @(posedge clk) begin
         op_in_2_21 <= op_out_2_20;
         pivot_in_2_21 <= pivot_out_2_20;
         start_in_2_21 <= start_out_2_20;
         swap_in_2_21 <= swap_out_2_20;
     end

     always @(posedge clk) begin
         data_in_2_21 <= data_out_1_21;
     end
  
     processor_AB AB_2_21 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_21),
       .start_in   (start_in_2_21),
       .swap_in   (swap_in_2_21),
       .op_in      (op_in_2_21),
       .pivot_in   (pivot_in_2_21),
       .start_out  (start_out_2_21),
       .swap_out   (swap_out_2_21),
       .data_out   (data_out_2_21),
       .op_out     (op_out_2_21),
       .pivot_out  (pivot_out_2_21),
       .r          (r_2_21)
     );

  // row 2, col 22

     reg start_in_2_22;
     wire start_out_2_22;

     reg swap_in_2_22;
     wire swap_out_2_22;

     reg [1:0] op_in_2_22;
     wire [1:0] op_out_2_22;

     wire r_2_22;

     reg data_in_2_22;
     wire data_out_2_22;

     reg pivot_in_2_22;
     wire pivot_out_2_22;

     always @(posedge clk) begin
         op_in_2_22 <= op_out_2_21;
         pivot_in_2_22 <= pivot_out_2_21;
         start_in_2_22 <= start_out_2_21;
         swap_in_2_22 <= swap_out_2_21;
     end

     always @(posedge clk) begin
         data_in_2_22 <= data_out_1_22;
     end
  
     processor_AB AB_2_22 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_22),
       .start_in   (start_in_2_22),
       .swap_in   (swap_in_2_22),
       .op_in      (op_in_2_22),
       .pivot_in   (pivot_in_2_22),
       .start_out  (start_out_2_22),
       .swap_out   (swap_out_2_22),
       .data_out   (data_out_2_22),
       .op_out     (op_out_2_22),
       .pivot_out  (pivot_out_2_22),
       .r          (r_2_22)
     );

  // row 2, col 23

     reg start_in_2_23;
     wire start_out_2_23;

     reg swap_in_2_23;
     wire swap_out_2_23;

     reg [1:0] op_in_2_23;
     wire [1:0] op_out_2_23;

     wire r_2_23;

     reg data_in_2_23;
     wire data_out_2_23;

     reg pivot_in_2_23;
     wire pivot_out_2_23;

     always @(posedge clk) begin
         op_in_2_23 <= op_out_2_22;
         pivot_in_2_23 <= pivot_out_2_22;
         start_in_2_23 <= start_out_2_22;
         swap_in_2_23 <= swap_out_2_22;
     end

     always @(posedge clk) begin
         data_in_2_23 <= data_out_1_23;
     end
  
     processor_AB AB_2_23 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_23),
       .start_in   (start_in_2_23),
       .swap_in   (swap_in_2_23),
       .op_in      (op_in_2_23),
       .pivot_in   (pivot_in_2_23),
       .start_out  (start_out_2_23),
       .swap_out   (swap_out_2_23),
       .data_out   (data_out_2_23),
       .op_out     (op_out_2_23),
       .pivot_out  (pivot_out_2_23),
       .r          (r_2_23)
     );

  // row 2, col 24

     reg start_in_2_24;
     wire start_out_2_24;

     reg swap_in_2_24;
     wire swap_out_2_24;

     reg [1:0] op_in_2_24;
     wire [1:0] op_out_2_24;

     wire r_2_24;

     reg data_in_2_24;
     wire data_out_2_24;

     reg pivot_in_2_24;
     wire pivot_out_2_24;

     always @(posedge clk) begin
         op_in_2_24 <= op_out_2_23;
         pivot_in_2_24 <= pivot_out_2_23;
         start_in_2_24 <= start_out_2_23;
         swap_in_2_24 <= swap_out_2_23;
     end

     always @(posedge clk) begin
         data_in_2_24 <= data_out_1_24;
     end
  
     processor_AB AB_2_24 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_24),
       .start_in   (start_in_2_24),
       .swap_in   (swap_in_2_24),
       .op_in      (op_in_2_24),
       .pivot_in   (pivot_in_2_24),
       .start_out  (start_out_2_24),
       .swap_out   (swap_out_2_24),
       .data_out   (data_out_2_24),
       .op_out     (op_out_2_24),
       .pivot_out  (pivot_out_2_24),
       .r          (r_2_24)
     );

  // row 2, col 25

     reg start_in_2_25;
     wire start_out_2_25;

     reg swap_in_2_25;
     wire swap_out_2_25;

     reg [1:0] op_in_2_25;
     wire [1:0] op_out_2_25;

     wire r_2_25;

     reg data_in_2_25;
     wire data_out_2_25;

     reg pivot_in_2_25;
     wire pivot_out_2_25;

     always @(posedge clk) begin
         op_in_2_25 <= op_out_2_24;
         pivot_in_2_25 <= pivot_out_2_24;
         start_in_2_25 <= start_out_2_24;
         swap_in_2_25 <= swap_out_2_24;
     end

     always @(posedge clk) begin
         data_in_2_25 <= data_out_1_25;
     end
  
     processor_AB AB_2_25 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_25),
       .start_in   (start_in_2_25),
       .swap_in   (swap_in_2_25),
       .op_in      (op_in_2_25),
       .pivot_in   (pivot_in_2_25),
       .start_out  (start_out_2_25),
       .swap_out   (swap_out_2_25),
       .data_out   (data_out_2_25),
       .op_out     (op_out_2_25),
       .pivot_out  (pivot_out_2_25),
       .r          (r_2_25)
     );

  // row 2, col 26

     reg start_in_2_26;
     wire start_out_2_26;

     reg swap_in_2_26;
     wire swap_out_2_26;

     reg [1:0] op_in_2_26;
     wire [1:0] op_out_2_26;

     wire r_2_26;

     reg data_in_2_26;
     wire data_out_2_26;

     reg pivot_in_2_26;
     wire pivot_out_2_26;

     always @(posedge clk) begin
         op_in_2_26 <= op_out_2_25;
         pivot_in_2_26 <= pivot_out_2_25;
         start_in_2_26 <= start_out_2_25;
         swap_in_2_26 <= swap_out_2_25;
     end

     always @(posedge clk) begin
         data_in_2_26 <= data_out_1_26;
     end
  
     processor_AB AB_2_26 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_26),
       .start_in   (start_in_2_26),
       .swap_in   (swap_in_2_26),
       .op_in      (op_in_2_26),
       .pivot_in   (pivot_in_2_26),
       .start_out  (start_out_2_26),
       .swap_out   (swap_out_2_26),
       .data_out   (data_out_2_26),
       .op_out     (op_out_2_26),
       .pivot_out  (pivot_out_2_26),
       .r          (r_2_26)
     );

  // row 2, col 27

     reg start_in_2_27;
     wire start_out_2_27;

     reg swap_in_2_27;
     wire swap_out_2_27;

     reg [1:0] op_in_2_27;
     wire [1:0] op_out_2_27;

     wire r_2_27;

     reg data_in_2_27;
     wire data_out_2_27;

     reg pivot_in_2_27;
     wire pivot_out_2_27;

     always @(posedge clk) begin
         op_in_2_27 <= op_out_2_26;
         pivot_in_2_27 <= pivot_out_2_26;
         start_in_2_27 <= start_out_2_26;
         swap_in_2_27 <= swap_out_2_26;
     end

     always @(posedge clk) begin
         data_in_2_27 <= data_out_1_27;
     end
  
     processor_AB AB_2_27 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_27),
       .start_in   (start_in_2_27),
       .swap_in   (swap_in_2_27),
       .op_in      (op_in_2_27),
       .pivot_in   (pivot_in_2_27),
       .start_out  (start_out_2_27),
       .swap_out   (swap_out_2_27),
       .data_out   (data_out_2_27),
       .op_out     (op_out_2_27),
       .pivot_out  (pivot_out_2_27),
       .r          (r_2_27)
     );

  // row 2, col 28

     reg start_in_2_28;
     wire start_out_2_28;

     reg swap_in_2_28;
     wire swap_out_2_28;

     reg [1:0] op_in_2_28;
     wire [1:0] op_out_2_28;

     wire r_2_28;

     reg data_in_2_28;
     wire data_out_2_28;

     reg pivot_in_2_28;
     wire pivot_out_2_28;

     always @(posedge clk) begin
         op_in_2_28 <= op_out_2_27;
         pivot_in_2_28 <= pivot_out_2_27;
         start_in_2_28 <= start_out_2_27;
         swap_in_2_28 <= swap_out_2_27;
     end

     always @(posedge clk) begin
         data_in_2_28 <= data_out_1_28;
     end
  
     processor_AB AB_2_28 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_28),
       .start_in   (start_in_2_28),
       .swap_in   (swap_in_2_28),
       .op_in      (op_in_2_28),
       .pivot_in   (pivot_in_2_28),
       .start_out  (start_out_2_28),
       .swap_out   (swap_out_2_28),
       .data_out   (data_out_2_28),
       .op_out     (op_out_2_28),
       .pivot_out  (pivot_out_2_28),
       .r          (r_2_28)
     );

  // row 2, col 29

     reg start_in_2_29;
     wire start_out_2_29;

     reg swap_in_2_29;
     wire swap_out_2_29;

     reg [1:0] op_in_2_29;
     wire [1:0] op_out_2_29;

     wire r_2_29;

     reg data_in_2_29;
     wire data_out_2_29;

     reg pivot_in_2_29;
     wire pivot_out_2_29;

     always @(posedge clk) begin
         op_in_2_29 <= op_out_2_28;
         pivot_in_2_29 <= pivot_out_2_28;
         start_in_2_29 <= start_out_2_28;
         swap_in_2_29 <= swap_out_2_28;
     end

     always @(posedge clk) begin
         data_in_2_29 <= data_out_1_29;
     end
  
     processor_AB AB_2_29 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_29),
       .start_in   (start_in_2_29),
       .swap_in   (swap_in_2_29),
       .op_in      (op_in_2_29),
       .pivot_in   (pivot_in_2_29),
       .start_out  (start_out_2_29),
       .swap_out   (swap_out_2_29),
       .data_out   (data_out_2_29),
       .op_out     (op_out_2_29),
       .pivot_out  (pivot_out_2_29),
       .r          (r_2_29)
     );

  // row 2, col 30

     reg start_in_2_30;
     wire start_out_2_30;

     reg swap_in_2_30;
     wire swap_out_2_30;

     reg [1:0] op_in_2_30;
     wire [1:0] op_out_2_30;

     wire r_2_30;

     reg data_in_2_30;
     wire data_out_2_30;

     reg pivot_in_2_30;
     wire pivot_out_2_30;

     always @(posedge clk) begin
         op_in_2_30 <= op_out_2_29;
         pivot_in_2_30 <= pivot_out_2_29;
         start_in_2_30 <= start_out_2_29;
         swap_in_2_30 <= swap_out_2_29;
     end

     always @(posedge clk) begin
         data_in_2_30 <= data_out_1_30;
     end
  
     processor_AB AB_2_30 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_30),
       .start_in   (start_in_2_30),
       .swap_in   (swap_in_2_30),
       .op_in      (op_in_2_30),
       .pivot_in   (pivot_in_2_30),
       .start_out  (start_out_2_30),
       .swap_out   (swap_out_2_30),
       .data_out   (data_out_2_30),
       .op_out     (op_out_2_30),
       .pivot_out  (pivot_out_2_30),
       .r          (r_2_30)
     );

  // row 2, col 31

     reg start_in_2_31;
     wire start_out_2_31;

     reg swap_in_2_31;
     wire swap_out_2_31;

     reg [1:0] op_in_2_31;
     wire [1:0] op_out_2_31;

     wire r_2_31;

     reg data_in_2_31;
     wire data_out_2_31;

     reg pivot_in_2_31;
     wire pivot_out_2_31;

     always @(posedge clk) begin
         op_in_2_31 <= op_out_2_30;
         pivot_in_2_31 <= pivot_out_2_30;
         start_in_2_31 <= start_out_2_30;
         swap_in_2_31 <= swap_out_2_30;
     end

     always @(posedge clk) begin
         data_in_2_31 <= data_out_1_31;
     end
  
     processor_AB AB_2_31 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_31),
       .start_in   (start_in_2_31),
       .swap_in   (swap_in_2_31),
       .op_in      (op_in_2_31),
       .pivot_in   (pivot_in_2_31),
       .start_out  (start_out_2_31),
       .swap_out   (swap_out_2_31),
       .data_out   (data_out_2_31),
       .op_out     (op_out_2_31),
       .pivot_out  (pivot_out_2_31),
       .r          (r_2_31)
     );

  // row 2, col 32

     reg start_in_2_32;
     wire start_out_2_32;

     reg swap_in_2_32;
     wire swap_out_2_32;

     reg [1:0] op_in_2_32;
     wire [1:0] op_out_2_32;

     wire r_2_32;

     reg data_in_2_32;
     wire data_out_2_32;

     reg pivot_in_2_32;
     wire pivot_out_2_32;

     always @(posedge clk) begin
         op_in_2_32 <= op_out_2_31;
         pivot_in_2_32 <= pivot_out_2_31;
         start_in_2_32 <= start_out_2_31;
         swap_in_2_32 <= swap_out_2_31;
     end

     always @(posedge clk) begin
         data_in_2_32 <= data_out_1_32;
     end
  
     processor_AB AB_2_32 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_32),
       .start_in   (start_in_2_32),
       .swap_in   (swap_in_2_32),
       .op_in      (op_in_2_32),
       .pivot_in   (pivot_in_2_32),
       .start_out  (start_out_2_32),
       .swap_out   (swap_out_2_32),
       .data_out   (data_out_2_32),
       .op_out     (op_out_2_32),
       .pivot_out  (pivot_out_2_32),
       .r          (r_2_32)
     );

  // row 2, col 33

     reg start_in_2_33;
     wire start_out_2_33;

     reg swap_in_2_33;
     wire swap_out_2_33;

     reg [1:0] op_in_2_33;
     wire [1:0] op_out_2_33;

     wire r_2_33;

     reg data_in_2_33;
     wire data_out_2_33;

     reg pivot_in_2_33;
     wire pivot_out_2_33;

     always @(posedge clk) begin
         op_in_2_33 <= op_out_2_32;
         pivot_in_2_33 <= pivot_out_2_32;
         start_in_2_33 <= start_out_2_32;
         swap_in_2_33 <= swap_out_2_32;
     end

     always @(posedge clk) begin
         data_in_2_33 <= data_out_1_33;
     end
  
     processor_AB AB_2_33 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_33),
       .start_in   (start_in_2_33),
       .swap_in   (swap_in_2_33),
       .op_in      (op_in_2_33),
       .pivot_in   (pivot_in_2_33),
       .start_out  (start_out_2_33),
       .swap_out   (swap_out_2_33),
       .data_out   (data_out_2_33),
       .op_out     (op_out_2_33),
       .pivot_out  (pivot_out_2_33),
       .r          (r_2_33)
     );

  // row 2, col 34

     reg start_in_2_34;
     wire start_out_2_34;

     reg swap_in_2_34;
     wire swap_out_2_34;

     reg [1:0] op_in_2_34;
     wire [1:0] op_out_2_34;

     wire r_2_34;

     reg data_in_2_34;
     wire data_out_2_34;

     reg pivot_in_2_34;
     wire pivot_out_2_34;

     always @(posedge clk) begin
         op_in_2_34 <= op_out_2_33;
         pivot_in_2_34 <= pivot_out_2_33;
         start_in_2_34 <= start_out_2_33;
         swap_in_2_34 <= swap_out_2_33;
     end

     always @(posedge clk) begin
         data_in_2_34 <= data_out_1_34;
     end
  
     processor_AB AB_2_34 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_34),
       .start_in   (start_in_2_34),
       .swap_in   (swap_in_2_34),
       .op_in      (op_in_2_34),
       .pivot_in   (pivot_in_2_34),
       .start_out  (start_out_2_34),
       .swap_out   (swap_out_2_34),
       .data_out   (data_out_2_34),
       .op_out     (op_out_2_34),
       .pivot_out  (pivot_out_2_34),
       .r          (r_2_34)
     );

  // row 2, col 35

     reg start_in_2_35;
     wire start_out_2_35;

     reg swap_in_2_35;
     wire swap_out_2_35;

     reg [1:0] op_in_2_35;
     wire [1:0] op_out_2_35;

     wire r_2_35;

     reg data_in_2_35;
     wire data_out_2_35;

     reg pivot_in_2_35;
     wire pivot_out_2_35;

     always @(posedge clk) begin
         op_in_2_35 <= op_out_2_34;
         pivot_in_2_35 <= pivot_out_2_34;
         start_in_2_35 <= start_out_2_34;
         swap_in_2_35 <= swap_out_2_34;
     end

     always @(posedge clk) begin
         data_in_2_35 <= data_out_1_35;
     end
  
     processor_AB AB_2_35 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_35),
       .start_in   (start_in_2_35),
       .swap_in   (swap_in_2_35),
       .op_in      (op_in_2_35),
       .pivot_in   (pivot_in_2_35),
       .start_out  (start_out_2_35),
       .swap_out   (swap_out_2_35),
       .data_out   (data_out_2_35),
       .op_out     (op_out_2_35),
       .pivot_out  (pivot_out_2_35),
       .r          (r_2_35)
     );

  // row 2, col 36

     reg start_in_2_36;
     wire start_out_2_36;

     reg swap_in_2_36;
     wire swap_out_2_36;

     reg [1:0] op_in_2_36;
     wire [1:0] op_out_2_36;

     wire r_2_36;

     reg data_in_2_36;
     wire data_out_2_36;

     reg pivot_in_2_36;
     wire pivot_out_2_36;

     always @(posedge clk) begin
         op_in_2_36 <= op_out_2_35;
         pivot_in_2_36 <= pivot_out_2_35;
         start_in_2_36 <= start_out_2_35;
         swap_in_2_36 <= swap_out_2_35;
     end

     always @(posedge clk) begin
         data_in_2_36 <= data_out_1_36;
     end
  
     processor_AB AB_2_36 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_36),
       .start_in   (start_in_2_36),
       .swap_in   (swap_in_2_36),
       .op_in      (op_in_2_36),
       .pivot_in   (pivot_in_2_36),
       .start_out  (start_out_2_36),
       .swap_out   (swap_out_2_36),
       .data_out   (data_out_2_36),
       .op_out     (op_out_2_36),
       .pivot_out  (pivot_out_2_36),
       .r          (r_2_36)
     );

  // row 2, col 37

     reg start_in_2_37;
     wire start_out_2_37;

     reg swap_in_2_37;
     wire swap_out_2_37;

     reg [1:0] op_in_2_37;
     wire [1:0] op_out_2_37;

     wire r_2_37;

     reg data_in_2_37;
     wire data_out_2_37;

     reg pivot_in_2_37;
     wire pivot_out_2_37;

     always @(posedge clk) begin
         op_in_2_37 <= op_out_2_36;
         pivot_in_2_37 <= pivot_out_2_36;
         start_in_2_37 <= start_out_2_36;
         swap_in_2_37 <= swap_out_2_36;
     end

     always @(posedge clk) begin
         data_in_2_37 <= data_out_1_37;
     end
  
     processor_AB AB_2_37 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_37),
       .start_in   (start_in_2_37),
       .swap_in   (swap_in_2_37),
       .op_in      (op_in_2_37),
       .pivot_in   (pivot_in_2_37),
       .start_out  (start_out_2_37),
       .swap_out   (swap_out_2_37),
       .data_out   (data_out_2_37),
       .op_out     (op_out_2_37),
       .pivot_out  (pivot_out_2_37),
       .r          (r_2_37)
     );

  // row 2, col 38

     reg start_in_2_38;
     wire start_out_2_38;

     reg swap_in_2_38;
     wire swap_out_2_38;

     reg [1:0] op_in_2_38;
     wire [1:0] op_out_2_38;

     wire r_2_38;

     reg data_in_2_38;
     wire data_out_2_38;

     reg pivot_in_2_38;
     wire pivot_out_2_38;

     always @(posedge clk) begin
         op_in_2_38 <= op_out_2_37;
         pivot_in_2_38 <= pivot_out_2_37;
         start_in_2_38 <= start_out_2_37;
         swap_in_2_38 <= swap_out_2_37;
     end

     always @(posedge clk) begin
         data_in_2_38 <= data_out_1_38;
     end
  
     processor_AB AB_2_38 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_38),
       .start_in   (start_in_2_38),
       .swap_in   (swap_in_2_38),
       .op_in      (op_in_2_38),
       .pivot_in   (pivot_in_2_38),
       .start_out  (start_out_2_38),
       .swap_out   (swap_out_2_38),
       .data_out   (data_out_2_38),
       .op_out     (op_out_2_38),
       .pivot_out  (pivot_out_2_38),
       .r          (r_2_38)
     );

  // row 2, col 39

     reg start_in_2_39;
     wire start_out_2_39;

     reg swap_in_2_39;
     wire swap_out_2_39;

     reg [1:0] op_in_2_39;
     wire [1:0] op_out_2_39;

     wire r_2_39;

     reg data_in_2_39;
     wire data_out_2_39;

     reg pivot_in_2_39;
     wire pivot_out_2_39;

     always @(posedge clk) begin
         op_in_2_39 <= op_out_2_38;
         pivot_in_2_39 <= pivot_out_2_38;
         start_in_2_39 <= start_out_2_38;
         swap_in_2_39 <= swap_out_2_38;
     end

     always @(posedge clk) begin
         data_in_2_39 <= data_out_1_39;
     end
  
     processor_AB AB_2_39 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_39),
       .start_in   (start_in_2_39),
       .swap_in   (swap_in_2_39),
       .op_in      (op_in_2_39),
       .pivot_in   (pivot_in_2_39),
       .start_out  (start_out_2_39),
       .swap_out   (swap_out_2_39),
       .data_out   (data_out_2_39),
       .op_out     (op_out_2_39),
       .pivot_out  (pivot_out_2_39),
       .r          (r_2_39)
     );

  // row 2, col 40

     reg start_in_2_40;
     wire start_out_2_40;

     reg swap_in_2_40;
     wire swap_out_2_40;

     reg [1:0] op_in_2_40;
     wire [1:0] op_out_2_40;

     wire r_2_40;

     reg data_in_2_40;
     wire data_out_2_40;

     reg pivot_in_2_40;
     wire pivot_out_2_40;

     always @(posedge clk) begin
         op_in_2_40 <= op_out_2_39;
         pivot_in_2_40 <= pivot_out_2_39;
         start_in_2_40 <= start_out_2_39;
         swap_in_2_40 <= swap_out_2_39;
     end

     always @(posedge clk) begin
         data_in_2_40 <= data_out_1_40;
     end
  
     processor_AB AB_2_40 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_40),
       .start_in   (start_in_2_40),
       .swap_in   (swap_in_2_40),
       .op_in      (op_in_2_40),
       .pivot_in   (pivot_in_2_40),
       .start_out  (start_out_2_40),
       .swap_out   (swap_out_2_40),
       .data_out   (data_out_2_40),
       .op_out     (op_out_2_40),
       .pivot_out  (pivot_out_2_40),
       .r          (r_2_40)
     );

  // row 2, col 41

     reg start_in_2_41;
     wire start_out_2_41;

     reg swap_in_2_41;
     wire swap_out_2_41;

     reg [1:0] op_in_2_41;
     wire [1:0] op_out_2_41;

     wire r_2_41;

     reg data_in_2_41;
     wire data_out_2_41;

     reg pivot_in_2_41;
     wire pivot_out_2_41;

     always @(posedge clk) begin
         op_in_2_41 <= op_out_2_40;
         pivot_in_2_41 <= pivot_out_2_40;
         start_in_2_41 <= start_out_2_40;
         swap_in_2_41 <= swap_out_2_40;
     end

     always @(posedge clk) begin
         data_in_2_41 <= data_out_1_41;
     end
  
     processor_AB AB_2_41 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_41),
       .start_in   (start_in_2_41),
       .swap_in   (swap_in_2_41),
       .op_in      (op_in_2_41),
       .pivot_in   (pivot_in_2_41),
       .start_out  (start_out_2_41),
       .swap_out   (swap_out_2_41),
       .data_out   (data_out_2_41),
       .op_out     (op_out_2_41),
       .pivot_out  (pivot_out_2_41),
       .r          (r_2_41)
     );

  // row 2, col 42

     reg start_in_2_42;
     wire start_out_2_42;

     reg swap_in_2_42;
     wire swap_out_2_42;

     reg [1:0] op_in_2_42;
     wire [1:0] op_out_2_42;

     wire r_2_42;

     reg data_in_2_42;
     wire data_out_2_42;

     reg pivot_in_2_42;
     wire pivot_out_2_42;

     always @(posedge clk) begin
         op_in_2_42 <= op_out_2_41;
         pivot_in_2_42 <= pivot_out_2_41;
         start_in_2_42 <= start_out_2_41;
         swap_in_2_42 <= swap_out_2_41;
     end

     always @(posedge clk) begin
         data_in_2_42 <= data_out_1_42;
     end
  
     processor_AB AB_2_42 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_42),
       .start_in   (start_in_2_42),
       .swap_in   (swap_in_2_42),
       .op_in      (op_in_2_42),
       .pivot_in   (pivot_in_2_42),
       .start_out  (start_out_2_42),
       .swap_out   (swap_out_2_42),
       .data_out   (data_out_2_42),
       .op_out     (op_out_2_42),
       .pivot_out  (pivot_out_2_42),
       .r          (r_2_42)
     );

  // row 2, col 43

     reg start_in_2_43;
     wire start_out_2_43;

     reg swap_in_2_43;
     wire swap_out_2_43;

     reg [1:0] op_in_2_43;
     wire [1:0] op_out_2_43;

     wire r_2_43;

     reg data_in_2_43;
     wire data_out_2_43;

     reg pivot_in_2_43;
     wire pivot_out_2_43;

     always @(posedge clk) begin
         op_in_2_43 <= op_out_2_42;
         pivot_in_2_43 <= pivot_out_2_42;
         start_in_2_43 <= start_out_2_42;
         swap_in_2_43 <= swap_out_2_42;
     end

     always @(posedge clk) begin
         data_in_2_43 <= data_out_1_43;
     end
  
     processor_AB AB_2_43 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_43),
       .start_in   (start_in_2_43),
       .swap_in   (swap_in_2_43),
       .op_in      (op_in_2_43),
       .pivot_in   (pivot_in_2_43),
       .start_out  (start_out_2_43),
       .swap_out   (swap_out_2_43),
       .data_out   (data_out_2_43),
       .op_out     (op_out_2_43),
       .pivot_out  (pivot_out_2_43),
       .r          (r_2_43)
     );

  // row 2, col 44

     reg start_in_2_44;
     wire start_out_2_44;

     reg swap_in_2_44;
     wire swap_out_2_44;

     reg [1:0] op_in_2_44;
     wire [1:0] op_out_2_44;

     wire r_2_44;

     reg data_in_2_44;
     wire data_out_2_44;

     reg pivot_in_2_44;
     wire pivot_out_2_44;

     always @(posedge clk) begin
         op_in_2_44 <= op_out_2_43;
         pivot_in_2_44 <= pivot_out_2_43;
         start_in_2_44 <= start_out_2_43;
         swap_in_2_44 <= swap_out_2_43;
     end

     always @(posedge clk) begin
         data_in_2_44 <= data_out_1_44;
     end
  
     processor_AB AB_2_44 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_44),
       .start_in   (start_in_2_44),
       .swap_in   (swap_in_2_44),
       .op_in      (op_in_2_44),
       .pivot_in   (pivot_in_2_44),
       .start_out  (start_out_2_44),
       .swap_out   (swap_out_2_44),
       .data_out   (data_out_2_44),
       .op_out     (op_out_2_44),
       .pivot_out  (pivot_out_2_44),
       .r          (r_2_44)
     );

  // row 2, col 45

     reg start_in_2_45;
     wire start_out_2_45;

     reg swap_in_2_45;
     wire swap_out_2_45;

     reg [1:0] op_in_2_45;
     wire [1:0] op_out_2_45;

     wire r_2_45;

     reg data_in_2_45;
     wire data_out_2_45;

     reg pivot_in_2_45;
     wire pivot_out_2_45;

     always @(posedge clk) begin
         op_in_2_45 <= op_out_2_44;
         pivot_in_2_45 <= pivot_out_2_44;
         start_in_2_45 <= start_out_2_44;
         swap_in_2_45 <= swap_out_2_44;
     end

     always @(posedge clk) begin
         data_in_2_45 <= data_out_1_45;
     end
  
     processor_AB AB_2_45 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_45),
       .start_in   (start_in_2_45),
       .swap_in   (swap_in_2_45),
       .op_in      (op_in_2_45),
       .pivot_in   (pivot_in_2_45),
       .start_out  (start_out_2_45),
       .swap_out   (swap_out_2_45),
       .data_out   (data_out_2_45),
       .op_out     (op_out_2_45),
       .pivot_out  (pivot_out_2_45),
       .r          (r_2_45)
     );

  // row 2, col 46

     reg start_in_2_46;
     wire start_out_2_46;

     reg swap_in_2_46;
     wire swap_out_2_46;

     reg [1:0] op_in_2_46;
     wire [1:0] op_out_2_46;

     wire r_2_46;

     reg data_in_2_46;
     wire data_out_2_46;

     reg pivot_in_2_46;
     wire pivot_out_2_46;

     always @(posedge clk) begin
         op_in_2_46 <= op_out_2_45;
         pivot_in_2_46 <= pivot_out_2_45;
         start_in_2_46 <= start_out_2_45;
         swap_in_2_46 <= swap_out_2_45;
     end

     always @(posedge clk) begin
         data_in_2_46 <= data_out_1_46;
     end
  
     processor_AB AB_2_46 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_46),
       .start_in   (start_in_2_46),
       .swap_in   (swap_in_2_46),
       .op_in      (op_in_2_46),
       .pivot_in   (pivot_in_2_46),
       .start_out  (start_out_2_46),
       .swap_out   (swap_out_2_46),
       .data_out   (data_out_2_46),
       .op_out     (op_out_2_46),
       .pivot_out  (pivot_out_2_46),
       .r          (r_2_46)
     );

  // row 2, col 47

     reg start_in_2_47;
     wire start_out_2_47;

     reg swap_in_2_47;
     wire swap_out_2_47;

     reg [1:0] op_in_2_47;
     wire [1:0] op_out_2_47;

     wire r_2_47;

     reg data_in_2_47;
     wire data_out_2_47;

     reg pivot_in_2_47;
     wire pivot_out_2_47;

     always @(posedge clk) begin
         op_in_2_47 <= op_out_2_46;
         pivot_in_2_47 <= pivot_out_2_46;
         start_in_2_47 <= start_out_2_46;
         swap_in_2_47 <= swap_out_2_46;
     end

     always @(posedge clk) begin
         data_in_2_47 <= data_out_1_47;
     end
  
     processor_AB AB_2_47 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_47),
       .start_in   (start_in_2_47),
       .swap_in   (swap_in_2_47),
       .op_in      (op_in_2_47),
       .pivot_in   (pivot_in_2_47),
       .start_out  (start_out_2_47),
       .swap_out   (swap_out_2_47),
       .data_out   (data_out_2_47),
       .op_out     (op_out_2_47),
       .pivot_out  (pivot_out_2_47),
       .r          (r_2_47)
     );

  // row 2, col 48

     reg start_in_2_48;
     wire start_out_2_48;

     reg swap_in_2_48;
     wire swap_out_2_48;

     reg [1:0] op_in_2_48;
     wire [1:0] op_out_2_48;

     wire r_2_48;

     reg data_in_2_48;
     wire data_out_2_48;

     reg pivot_in_2_48;
     wire pivot_out_2_48;

     always @(posedge clk) begin
         op_in_2_48 <= op_out_2_47;
         pivot_in_2_48 <= pivot_out_2_47;
         start_in_2_48 <= start_out_2_47;
         swap_in_2_48 <= swap_out_2_47;
     end

     always @(posedge clk) begin
         data_in_2_48 <= data_out_1_48;
     end
  
     processor_AB AB_2_48 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_48),
       .start_in   (start_in_2_48),
       .swap_in   (swap_in_2_48),
       .op_in      (op_in_2_48),
       .pivot_in   (pivot_in_2_48),
       .start_out  (start_out_2_48),
       .swap_out   (swap_out_2_48),
       .data_out   (data_out_2_48),
       .op_out     (op_out_2_48),
       .pivot_out  (pivot_out_2_48),
       .r          (r_2_48)
     );

  // row 2, col 49

     reg start_in_2_49;
     wire start_out_2_49;

     reg swap_in_2_49;
     wire swap_out_2_49;

     reg [1:0] op_in_2_49;
     wire [1:0] op_out_2_49;

     wire r_2_49;

     reg data_in_2_49;
     wire data_out_2_49;

     reg pivot_in_2_49;
     wire pivot_out_2_49;

     always @(posedge clk) begin
         op_in_2_49 <= op_out_2_48;
         pivot_in_2_49 <= pivot_out_2_48;
         start_in_2_49 <= start_out_2_48;
         swap_in_2_49 <= swap_out_2_48;
     end

     always @(posedge clk) begin
         data_in_2_49 <= data_out_1_49;
     end
  
     processor_AB AB_2_49 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_49),
       .start_in   (start_in_2_49),
       .swap_in   (swap_in_2_49),
       .op_in      (op_in_2_49),
       .pivot_in   (pivot_in_2_49),
       .start_out  (start_out_2_49),
       .swap_out   (swap_out_2_49),
       .data_out   (data_out_2_49),
       .op_out     (op_out_2_49),
       .pivot_out  (pivot_out_2_49),
       .r          (r_2_49)
     );

  // row 2, col 50

     reg start_in_2_50;
     wire start_out_2_50;

     reg swap_in_2_50;
     wire swap_out_2_50;

     reg [1:0] op_in_2_50;
     wire [1:0] op_out_2_50;

     wire r_2_50;

     reg data_in_2_50;
     wire data_out_2_50;

     reg pivot_in_2_50;
     wire pivot_out_2_50;

     always @(posedge clk) begin
         op_in_2_50 <= op_out_2_49;
         pivot_in_2_50 <= pivot_out_2_49;
         start_in_2_50 <= start_out_2_49;
         swap_in_2_50 <= swap_out_2_49;
     end

     always @(posedge clk) begin
         data_in_2_50 <= data_out_1_50;
     end
  
     processor_AB AB_2_50 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_50),
       .start_in   (start_in_2_50),
       .swap_in   (swap_in_2_50),
       .op_in      (op_in_2_50),
       .pivot_in   (pivot_in_2_50),
       .start_out  (start_out_2_50),
       .swap_out   (swap_out_2_50),
       .data_out   (data_out_2_50),
       .op_out     (op_out_2_50),
       .pivot_out  (pivot_out_2_50),
       .r          (r_2_50)
     );

  // row 2, col 51

     reg start_in_2_51;
     wire start_out_2_51;

     reg swap_in_2_51;
     wire swap_out_2_51;

     reg [1:0] op_in_2_51;
     wire [1:0] op_out_2_51;

     wire r_2_51;

     reg data_in_2_51;
     wire data_out_2_51;

     reg pivot_in_2_51;
     wire pivot_out_2_51;

     always @(posedge clk) begin
         op_in_2_51 <= op_out_2_50;
         pivot_in_2_51 <= pivot_out_2_50;
         start_in_2_51 <= start_out_2_50;
         swap_in_2_51 <= swap_out_2_50;
     end

     always @(posedge clk) begin
         data_in_2_51 <= data_out_1_51;
     end
  
     processor_AB AB_2_51 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_51),
       .start_in   (start_in_2_51),
       .swap_in   (swap_in_2_51),
       .op_in      (op_in_2_51),
       .pivot_in   (pivot_in_2_51),
       .start_out  (start_out_2_51),
       .swap_out   (swap_out_2_51),
       .data_out   (data_out_2_51),
       .op_out     (op_out_2_51),
       .pivot_out  (pivot_out_2_51),
       .r          (r_2_51)
     );

  // row 2, col 52

     reg start_in_2_52;
     wire start_out_2_52;

     reg swap_in_2_52;
     wire swap_out_2_52;

     reg [1:0] op_in_2_52;
     wire [1:0] op_out_2_52;

     wire r_2_52;

     reg data_in_2_52;
     wire data_out_2_52;

     reg pivot_in_2_52;
     wire pivot_out_2_52;

     always @(posedge clk) begin
         op_in_2_52 <= op_out_2_51;
         pivot_in_2_52 <= pivot_out_2_51;
         start_in_2_52 <= start_out_2_51;
         swap_in_2_52 <= swap_out_2_51;
     end

     always @(posedge clk) begin
         data_in_2_52 <= data_out_1_52;
     end
  
     processor_AB AB_2_52 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_52),
       .start_in   (start_in_2_52),
       .swap_in   (swap_in_2_52),
       .op_in      (op_in_2_52),
       .pivot_in   (pivot_in_2_52),
       .start_out  (start_out_2_52),
       .swap_out   (swap_out_2_52),
       .data_out   (data_out_2_52),
       .op_out     (op_out_2_52),
       .pivot_out  (pivot_out_2_52),
       .r          (r_2_52)
     );

  // row 2, col 53

     reg start_in_2_53;
     wire start_out_2_53;

     reg swap_in_2_53;
     wire swap_out_2_53;

     reg [1:0] op_in_2_53;
     wire [1:0] op_out_2_53;

     wire r_2_53;

     reg data_in_2_53;
     wire data_out_2_53;

     reg pivot_in_2_53;
     wire pivot_out_2_53;

     always @(posedge clk) begin
         op_in_2_53 <= op_out_2_52;
         pivot_in_2_53 <= pivot_out_2_52;
         start_in_2_53 <= start_out_2_52;
         swap_in_2_53 <= swap_out_2_52;
     end

     always @(posedge clk) begin
         data_in_2_53 <= data_out_1_53;
     end
  
     processor_AB AB_2_53 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_53),
       .start_in   (start_in_2_53),
       .swap_in   (swap_in_2_53),
       .op_in      (op_in_2_53),
       .pivot_in   (pivot_in_2_53),
       .start_out  (start_out_2_53),
       .swap_out   (swap_out_2_53),
       .data_out   (data_out_2_53),
       .op_out     (op_out_2_53),
       .pivot_out  (pivot_out_2_53),
       .r          (r_2_53)
     );

  // row 2, col 54

     reg start_in_2_54;
     wire start_out_2_54;

     reg swap_in_2_54;
     wire swap_out_2_54;

     reg [1:0] op_in_2_54;
     wire [1:0] op_out_2_54;

     wire r_2_54;

     reg data_in_2_54;
     wire data_out_2_54;

     reg pivot_in_2_54;
     wire pivot_out_2_54;

     always @(posedge clk) begin
         op_in_2_54 <= op_out_2_53;
         pivot_in_2_54 <= pivot_out_2_53;
         start_in_2_54 <= start_out_2_53;
         swap_in_2_54 <= swap_out_2_53;
     end

     always @(posedge clk) begin
         data_in_2_54 <= data_out_1_54;
     end
  
     processor_AB AB_2_54 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_54),
       .start_in   (start_in_2_54),
       .swap_in   (swap_in_2_54),
       .op_in      (op_in_2_54),
       .pivot_in   (pivot_in_2_54),
       .start_out  (start_out_2_54),
       .swap_out   (swap_out_2_54),
       .data_out   (data_out_2_54),
       .op_out     (op_out_2_54),
       .pivot_out  (pivot_out_2_54),
       .r          (r_2_54)
     );

  // row 2, col 55

     reg start_in_2_55;
     wire start_out_2_55;

     reg swap_in_2_55;
     wire swap_out_2_55;

     reg [1:0] op_in_2_55;
     wire [1:0] op_out_2_55;

     wire r_2_55;

     reg data_in_2_55;
     wire data_out_2_55;

     reg pivot_in_2_55;
     wire pivot_out_2_55;

     always @(posedge clk) begin
         op_in_2_55 <= op_out_2_54;
         pivot_in_2_55 <= pivot_out_2_54;
         start_in_2_55 <= start_out_2_54;
         swap_in_2_55 <= swap_out_2_54;
     end

     always @(posedge clk) begin
         data_in_2_55 <= data_out_1_55;
     end
  
     processor_AB AB_2_55 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_55),
       .start_in   (start_in_2_55),
       .swap_in   (swap_in_2_55),
       .op_in      (op_in_2_55),
       .pivot_in   (pivot_in_2_55),
       .start_out  (start_out_2_55),
       .swap_out   (swap_out_2_55),
       .data_out   (data_out_2_55),
       .op_out     (op_out_2_55),
       .pivot_out  (pivot_out_2_55),
       .r          (r_2_55)
     );

  // row 2, col 56

     reg start_in_2_56;
     wire start_out_2_56;

     reg swap_in_2_56;
     wire swap_out_2_56;

     reg [1:0] op_in_2_56;
     wire [1:0] op_out_2_56;

     wire r_2_56;

     reg data_in_2_56;
     wire data_out_2_56;

     reg pivot_in_2_56;
     wire pivot_out_2_56;

     always @(posedge clk) begin
         op_in_2_56 <= op_out_2_55;
         pivot_in_2_56 <= pivot_out_2_55;
         start_in_2_56 <= start_out_2_55;
         swap_in_2_56 <= swap_out_2_55;
     end

     always @(posedge clk) begin
         data_in_2_56 <= data_out_1_56;
     end
  
     processor_AB AB_2_56 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_56),
       .start_in   (start_in_2_56),
       .swap_in   (swap_in_2_56),
       .op_in      (op_in_2_56),
       .pivot_in   (pivot_in_2_56),
       .start_out  (start_out_2_56),
       .swap_out   (swap_out_2_56),
       .data_out   (data_out_2_56),
       .op_out     (op_out_2_56),
       .pivot_out  (pivot_out_2_56),
       .r          (r_2_56)
     );

  // row 2, col 57

     reg start_in_2_57;
     wire start_out_2_57;

     reg swap_in_2_57;
     wire swap_out_2_57;

     reg [1:0] op_in_2_57;
     wire [1:0] op_out_2_57;

     wire r_2_57;

     reg data_in_2_57;
     wire data_out_2_57;

     reg pivot_in_2_57;
     wire pivot_out_2_57;

     always @(posedge clk) begin
         op_in_2_57 <= op_out_2_56;
         pivot_in_2_57 <= pivot_out_2_56;
         start_in_2_57 <= start_out_2_56;
         swap_in_2_57 <= swap_out_2_56;
     end

     always @(posedge clk) begin
         data_in_2_57 <= data_out_1_57;
     end
  
     processor_AB AB_2_57 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_57),
       .start_in   (start_in_2_57),
       .swap_in   (swap_in_2_57),
       .op_in      (op_in_2_57),
       .pivot_in   (pivot_in_2_57),
       .start_out  (start_out_2_57),
       .swap_out   (swap_out_2_57),
       .data_out   (data_out_2_57),
       .op_out     (op_out_2_57),
       .pivot_out  (pivot_out_2_57),
       .r          (r_2_57)
     );

  // row 2, col 58

     reg start_in_2_58;
     wire start_out_2_58;

     reg swap_in_2_58;
     wire swap_out_2_58;

     reg [1:0] op_in_2_58;
     wire [1:0] op_out_2_58;

     wire r_2_58;

     reg data_in_2_58;
     wire data_out_2_58;

     reg pivot_in_2_58;
     wire pivot_out_2_58;

     always @(posedge clk) begin
         op_in_2_58 <= op_out_2_57;
         pivot_in_2_58 <= pivot_out_2_57;
         start_in_2_58 <= start_out_2_57;
         swap_in_2_58 <= swap_out_2_57;
     end

     always @(posedge clk) begin
         data_in_2_58 <= data_out_1_58;
     end
  
     processor_AB AB_2_58 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_58),
       .start_in   (start_in_2_58),
       .swap_in   (swap_in_2_58),
       .op_in      (op_in_2_58),
       .pivot_in   (pivot_in_2_58),
       .start_out  (start_out_2_58),
       .swap_out   (swap_out_2_58),
       .data_out   (data_out_2_58),
       .op_out     (op_out_2_58),
       .pivot_out  (pivot_out_2_58),
       .r          (r_2_58)
     );

  // row 2, col 59

     reg start_in_2_59;
     wire start_out_2_59;

     reg swap_in_2_59;
     wire swap_out_2_59;

     reg [1:0] op_in_2_59;
     wire [1:0] op_out_2_59;

     wire r_2_59;

     reg data_in_2_59;
     wire data_out_2_59;

     reg pivot_in_2_59;
     wire pivot_out_2_59;

     always @(posedge clk) begin
         op_in_2_59 <= op_out_2_58;
         pivot_in_2_59 <= pivot_out_2_58;
         start_in_2_59 <= start_out_2_58;
         swap_in_2_59 <= swap_out_2_58;
     end

     always @(posedge clk) begin
         data_in_2_59 <= data_out_1_59;
     end
  
     processor_AB AB_2_59 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_59),
       .start_in   (start_in_2_59),
       .swap_in   (swap_in_2_59),
       .op_in      (op_in_2_59),
       .pivot_in   (pivot_in_2_59),
       .start_out  (start_out_2_59),
       .swap_out   (swap_out_2_59),
       .data_out   (data_out_2_59),
       .op_out     (op_out_2_59),
       .pivot_out  (pivot_out_2_59),
       .r          (r_2_59)
     );

  // row 2, col 60

     reg start_in_2_60;
     wire start_out_2_60;

     reg swap_in_2_60;
     wire swap_out_2_60;

     reg [1:0] op_in_2_60;
     wire [1:0] op_out_2_60;

     wire r_2_60;

     reg data_in_2_60;
     wire data_out_2_60;

     reg pivot_in_2_60;
     wire pivot_out_2_60;

     always @(posedge clk) begin
         op_in_2_60 <= op_out_2_59;
         pivot_in_2_60 <= pivot_out_2_59;
         start_in_2_60 <= start_out_2_59;
         swap_in_2_60 <= swap_out_2_59;
     end

     always @(posedge clk) begin
         data_in_2_60 <= data_out_1_60;
     end
  
     processor_AB AB_2_60 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_60),
       .start_in   (start_in_2_60),
       .swap_in   (swap_in_2_60),
       .op_in      (op_in_2_60),
       .pivot_in   (pivot_in_2_60),
       .start_out  (start_out_2_60),
       .swap_out   (swap_out_2_60),
       .data_out   (data_out_2_60),
       .op_out     (op_out_2_60),
       .pivot_out  (pivot_out_2_60),
       .r          (r_2_60)
     );

  // row 2, col 61

     reg start_in_2_61;
     wire start_out_2_61;

     reg swap_in_2_61;
     wire swap_out_2_61;

     reg [1:0] op_in_2_61;
     wire [1:0] op_out_2_61;

     wire r_2_61;

     reg data_in_2_61;
     wire data_out_2_61;

     reg pivot_in_2_61;
     wire pivot_out_2_61;

     always @(posedge clk) begin
         op_in_2_61 <= op_out_2_60;
         pivot_in_2_61 <= pivot_out_2_60;
         start_in_2_61 <= start_out_2_60;
         swap_in_2_61 <= swap_out_2_60;
     end

     always @(posedge clk) begin
         data_in_2_61 <= data_out_1_61;
     end
  
     processor_AB AB_2_61 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_61),
       .start_in   (start_in_2_61),
       .swap_in   (swap_in_2_61),
       .op_in      (op_in_2_61),
       .pivot_in   (pivot_in_2_61),
       .start_out  (start_out_2_61),
       .swap_out   (swap_out_2_61),
       .data_out   (data_out_2_61),
       .op_out     (op_out_2_61),
       .pivot_out  (pivot_out_2_61),
       .r          (r_2_61)
     );

  // row 2, col 62

     reg start_in_2_62;
     wire start_out_2_62;

     reg swap_in_2_62;
     wire swap_out_2_62;

     reg [1:0] op_in_2_62;
     wire [1:0] op_out_2_62;

     wire r_2_62;

     reg data_in_2_62;
     wire data_out_2_62;

     reg pivot_in_2_62;
     wire pivot_out_2_62;

     always @(posedge clk) begin
         op_in_2_62 <= op_out_2_61;
         pivot_in_2_62 <= pivot_out_2_61;
         start_in_2_62 <= start_out_2_61;
         swap_in_2_62 <= swap_out_2_61;
     end

     always @(posedge clk) begin
         data_in_2_62 <= data_out_1_62;
     end
  
     processor_AB AB_2_62 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_62),
       .start_in   (start_in_2_62),
       .swap_in   (swap_in_2_62),
       .op_in      (op_in_2_62),
       .pivot_in   (pivot_in_2_62),
       .start_out  (start_out_2_62),
       .swap_out   (swap_out_2_62),
       .data_out   (data_out_2_62),
       .op_out     (op_out_2_62),
       .pivot_out  (pivot_out_2_62),
       .r          (r_2_62)
     );

  // row 2, col 63

     reg start_in_2_63;
     wire start_out_2_63;

     reg swap_in_2_63;
     wire swap_out_2_63;

     reg [1:0] op_in_2_63;
     wire [1:0] op_out_2_63;

     wire r_2_63;

     reg data_in_2_63;
     wire data_out_2_63;

     reg pivot_in_2_63;
     wire pivot_out_2_63;

     always @(posedge clk) begin
         op_in_2_63 <= op_out_2_62;
         pivot_in_2_63 <= pivot_out_2_62;
         start_in_2_63 <= start_out_2_62;
         swap_in_2_63 <= swap_out_2_62;
     end

     always @(posedge clk) begin
         data_in_2_63 <= data_out_1_63;
     end
  
     processor_AB AB_2_63 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_63),
       .start_in   (start_in_2_63),
       .swap_in   (swap_in_2_63),
       .op_in      (op_in_2_63),
       .pivot_in   (pivot_in_2_63),
       .start_out  (start_out_2_63),
       .swap_out   (swap_out_2_63),
       .data_out   (data_out_2_63),
       .op_out     (op_out_2_63),
       .pivot_out  (pivot_out_2_63),
       .r          (r_2_63)
     );

  // row 2, col 64

     reg start_in_2_64;
     wire start_out_2_64;

     reg swap_in_2_64;
     wire swap_out_2_64;

     reg [1:0] op_in_2_64;
     wire [1:0] op_out_2_64;

     wire r_2_64;

     reg data_in_2_64;
     wire data_out_2_64;

     reg pivot_in_2_64;
     wire pivot_out_2_64;

     always @(posedge clk) begin
         op_in_2_64 <= op_out_2_63;
         pivot_in_2_64 <= pivot_out_2_63;
         start_in_2_64 <= start_out_2_63;
         swap_in_2_64 <= swap_out_2_63;
     end

     always @(posedge clk) begin
         data_in_2_64 <= data_out_1_64;
     end
  
     processor_AB AB_2_64 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_64),
       .start_in   (start_in_2_64),
       .swap_in   (swap_in_2_64),
       .op_in      (op_in_2_64),
       .pivot_in   (pivot_in_2_64),
       .start_out  (start_out_2_64),
       .swap_out   (swap_out_2_64),
       .data_out   (data_out_2_64),
       .op_out     (op_out_2_64),
       .pivot_out  (pivot_out_2_64),
       .r          (r_2_64)
     );

  // row 2, col 65

     reg start_in_2_65;
     wire start_out_2_65;

     reg swap_in_2_65;
     wire swap_out_2_65;

     reg [1:0] op_in_2_65;
     wire [1:0] op_out_2_65;

     wire r_2_65;

     reg data_in_2_65;
     wire data_out_2_65;

     reg pivot_in_2_65;
     wire pivot_out_2_65;

     always @(posedge clk) begin
         op_in_2_65 <= op_out_2_64;
         pivot_in_2_65 <= pivot_out_2_64;
         start_in_2_65 <= start_out_2_64;
         swap_in_2_65 <= swap_out_2_64;
     end

     always @(posedge clk) begin
         data_in_2_65 <= data_out_1_65;
     end
  
     processor_AB AB_2_65 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_65),
       .start_in   (start_in_2_65),
       .swap_in   (swap_in_2_65),
       .op_in      (op_in_2_65),
       .pivot_in   (pivot_in_2_65),
       .start_out  (start_out_2_65),
       .swap_out   (swap_out_2_65),
       .data_out   (data_out_2_65),
       .op_out     (op_out_2_65),
       .pivot_out  (pivot_out_2_65),
       .r          (r_2_65)
     );

  // row 2, col 66

     reg start_in_2_66;
     wire start_out_2_66;

     reg swap_in_2_66;
     wire swap_out_2_66;

     reg [1:0] op_in_2_66;
     wire [1:0] op_out_2_66;

     wire r_2_66;

     reg data_in_2_66;
     wire data_out_2_66;

     reg pivot_in_2_66;
     wire pivot_out_2_66;

     always @(posedge clk) begin
         op_in_2_66 <= op_out_2_65;
         pivot_in_2_66 <= pivot_out_2_65;
         start_in_2_66 <= start_out_2_65;
         swap_in_2_66 <= swap_out_2_65;
     end

     always @(posedge clk) begin
         data_in_2_66 <= data_out_1_66;
     end
  
     processor_AB AB_2_66 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_66),
       .start_in   (start_in_2_66),
       .swap_in   (swap_in_2_66),
       .op_in      (op_in_2_66),
       .pivot_in   (pivot_in_2_66),
       .start_out  (start_out_2_66),
       .swap_out   (swap_out_2_66),
       .data_out   (data_out_2_66),
       .op_out     (op_out_2_66),
       .pivot_out  (pivot_out_2_66),
       .r          (r_2_66)
     );

  // row 2, col 67

     reg start_in_2_67;
     wire start_out_2_67;

     reg swap_in_2_67;
     wire swap_out_2_67;

     reg [1:0] op_in_2_67;
     wire [1:0] op_out_2_67;

     wire r_2_67;

     reg data_in_2_67;
     wire data_out_2_67;

     reg pivot_in_2_67;
     wire pivot_out_2_67;

     always @(posedge clk) begin
         op_in_2_67 <= op_out_2_66;
         pivot_in_2_67 <= pivot_out_2_66;
         start_in_2_67 <= start_out_2_66;
         swap_in_2_67 <= swap_out_2_66;
     end

     always @(posedge clk) begin
         data_in_2_67 <= data_out_1_67;
     end
  
     processor_AB AB_2_67 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_67),
       .start_in   (start_in_2_67),
       .swap_in   (swap_in_2_67),
       .op_in      (op_in_2_67),
       .pivot_in   (pivot_in_2_67),
       .start_out  (start_out_2_67),
       .swap_out   (swap_out_2_67),
       .data_out   (data_out_2_67),
       .op_out     (op_out_2_67),
       .pivot_out  (pivot_out_2_67),
       .r          (r_2_67)
     );

  // row 2, col 68

     reg start_in_2_68;
     wire start_out_2_68;

     reg swap_in_2_68;
     wire swap_out_2_68;

     reg [1:0] op_in_2_68;
     wire [1:0] op_out_2_68;

     wire r_2_68;

     reg data_in_2_68;
     wire data_out_2_68;

     reg pivot_in_2_68;
     wire pivot_out_2_68;

     always @(posedge clk) begin
         op_in_2_68 <= op_out_2_67;
         pivot_in_2_68 <= pivot_out_2_67;
         start_in_2_68 <= start_out_2_67;
         swap_in_2_68 <= swap_out_2_67;
     end

     always @(posedge clk) begin
         data_in_2_68 <= data_out_1_68;
     end
  
     processor_AB AB_2_68 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_68),
       .start_in   (start_in_2_68),
       .swap_in   (swap_in_2_68),
       .op_in      (op_in_2_68),
       .pivot_in   (pivot_in_2_68),
       .start_out  (start_out_2_68),
       .swap_out   (swap_out_2_68),
       .data_out   (data_out_2_68),
       .op_out     (op_out_2_68),
       .pivot_out  (pivot_out_2_68),
       .r          (r_2_68)
     );

  // row 2, col 69

     reg start_in_2_69;
     wire start_out_2_69;

     reg swap_in_2_69;
     wire swap_out_2_69;

     reg [1:0] op_in_2_69;
     wire [1:0] op_out_2_69;

     wire r_2_69;

     reg data_in_2_69;
     wire data_out_2_69;

     reg pivot_in_2_69;
     wire pivot_out_2_69;

     always @(posedge clk) begin
         op_in_2_69 <= op_out_2_68;
         pivot_in_2_69 <= pivot_out_2_68;
         start_in_2_69 <= start_out_2_68;
         swap_in_2_69 <= swap_out_2_68;
     end

     always @(posedge clk) begin
         data_in_2_69 <= data_out_1_69;
     end
  
     processor_AB AB_2_69 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_69),
       .start_in   (start_in_2_69),
       .swap_in   (swap_in_2_69),
       .op_in      (op_in_2_69),
       .pivot_in   (pivot_in_2_69),
       .start_out  (start_out_2_69),
       .swap_out   (swap_out_2_69),
       .data_out   (data_out_2_69),
       .op_out     (op_out_2_69),
       .pivot_out  (pivot_out_2_69),
       .r          (r_2_69)
     );

  // row 2, col 70

     reg start_in_2_70;
     wire start_out_2_70;

     reg swap_in_2_70;
     wire swap_out_2_70;

     reg [1:0] op_in_2_70;
     wire [1:0] op_out_2_70;

     wire r_2_70;

     reg data_in_2_70;
     wire data_out_2_70;

     reg pivot_in_2_70;
     wire pivot_out_2_70;

     always @(posedge clk) begin
         op_in_2_70 <= op_out_2_69;
         pivot_in_2_70 <= pivot_out_2_69;
         start_in_2_70 <= start_out_2_69;
         swap_in_2_70 <= swap_out_2_69;
     end

     always @(posedge clk) begin
         data_in_2_70 <= data_out_1_70;
     end
  
     processor_AB AB_2_70 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_70),
       .start_in   (start_in_2_70),
       .swap_in   (swap_in_2_70),
       .op_in      (op_in_2_70),
       .pivot_in   (pivot_in_2_70),
       .start_out  (start_out_2_70),
       .swap_out   (swap_out_2_70),
       .data_out   (data_out_2_70),
       .op_out     (op_out_2_70),
       .pivot_out  (pivot_out_2_70),
       .r          (r_2_70)
     );

  // row 2, col 71

     reg start_in_2_71;
     wire start_out_2_71;

     reg swap_in_2_71;
     wire swap_out_2_71;

     reg [1:0] op_in_2_71;
     wire [1:0] op_out_2_71;

     wire r_2_71;

     reg data_in_2_71;
     wire data_out_2_71;

     reg pivot_in_2_71;
     wire pivot_out_2_71;

     always @(posedge clk) begin
         op_in_2_71 <= op_out_2_70;
         pivot_in_2_71 <= pivot_out_2_70;
         start_in_2_71 <= start_out_2_70;
         swap_in_2_71 <= swap_out_2_70;
     end

     always @(posedge clk) begin
         data_in_2_71 <= data_out_1_71;
     end
  
     processor_AB AB_2_71 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_71),
       .start_in   (start_in_2_71),
       .swap_in   (swap_in_2_71),
       .op_in      (op_in_2_71),
       .pivot_in   (pivot_in_2_71),
       .start_out  (start_out_2_71),
       .swap_out   (swap_out_2_71),
       .data_out   (data_out_2_71),
       .op_out     (op_out_2_71),
       .pivot_out  (pivot_out_2_71),
       .r          (r_2_71)
     );

  // row 2, col 72

     reg start_in_2_72;
     wire start_out_2_72;

     reg swap_in_2_72;
     wire swap_out_2_72;

     reg [1:0] op_in_2_72;
     wire [1:0] op_out_2_72;

     wire r_2_72;

     reg data_in_2_72;
     wire data_out_2_72;

     reg pivot_in_2_72;
     wire pivot_out_2_72;

     always @(posedge clk) begin
         op_in_2_72 <= op_out_2_71;
         pivot_in_2_72 <= pivot_out_2_71;
         start_in_2_72 <= start_out_2_71;
         swap_in_2_72 <= swap_out_2_71;
     end

     always @(posedge clk) begin
         data_in_2_72 <= data_out_1_72;
     end
  
     processor_AB AB_2_72 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_72),
       .start_in   (start_in_2_72),
       .swap_in   (swap_in_2_72),
       .op_in      (op_in_2_72),
       .pivot_in   (pivot_in_2_72),
       .start_out  (start_out_2_72),
       .swap_out   (swap_out_2_72),
       .data_out   (data_out_2_72),
       .op_out     (op_out_2_72),
       .pivot_out  (pivot_out_2_72),
       .r          (r_2_72)
     );

  // row 2, col 73

     reg start_in_2_73;
     wire start_out_2_73;

     reg swap_in_2_73;
     wire swap_out_2_73;

     reg [1:0] op_in_2_73;
     wire [1:0] op_out_2_73;

     wire r_2_73;

     reg data_in_2_73;
     wire data_out_2_73;

     reg pivot_in_2_73;
     wire pivot_out_2_73;

     always @(posedge clk) begin
         op_in_2_73 <= op_out_2_72;
         pivot_in_2_73 <= pivot_out_2_72;
         start_in_2_73 <= start_out_2_72;
         swap_in_2_73 <= swap_out_2_72;
     end

     always @(posedge clk) begin
         data_in_2_73 <= data_out_1_73;
     end
  
     processor_AB AB_2_73 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_73),
       .start_in   (start_in_2_73),
       .swap_in   (swap_in_2_73),
       .op_in      (op_in_2_73),
       .pivot_in   (pivot_in_2_73),
       .start_out  (start_out_2_73),
       .swap_out   (swap_out_2_73),
       .data_out   (data_out_2_73),
       .op_out     (op_out_2_73),
       .pivot_out  (pivot_out_2_73),
       .r          (r_2_73)
     );

  // row 2, col 74

     reg start_in_2_74;
     wire start_out_2_74;

     reg swap_in_2_74;
     wire swap_out_2_74;

     reg [1:0] op_in_2_74;
     wire [1:0] op_out_2_74;

     wire r_2_74;

     reg data_in_2_74;
     wire data_out_2_74;

     reg pivot_in_2_74;
     wire pivot_out_2_74;

     always @(posedge clk) begin
         op_in_2_74 <= op_out_2_73;
         pivot_in_2_74 <= pivot_out_2_73;
         start_in_2_74 <= start_out_2_73;
         swap_in_2_74 <= swap_out_2_73;
     end

     always @(posedge clk) begin
         data_in_2_74 <= data_out_1_74;
     end
  
     processor_AB AB_2_74 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_74),
       .start_in   (start_in_2_74),
       .swap_in   (swap_in_2_74),
       .op_in      (op_in_2_74),
       .pivot_in   (pivot_in_2_74),
       .start_out  (start_out_2_74),
       .swap_out   (swap_out_2_74),
       .data_out   (data_out_2_74),
       .op_out     (op_out_2_74),
       .pivot_out  (pivot_out_2_74),
       .r          (r_2_74)
     );

  // row 2, col 75

     reg start_in_2_75;
     wire start_out_2_75;

     reg swap_in_2_75;
     wire swap_out_2_75;

     reg [1:0] op_in_2_75;
     wire [1:0] op_out_2_75;

     wire r_2_75;

     reg data_in_2_75;
     wire data_out_2_75;

     reg pivot_in_2_75;
     wire pivot_out_2_75;

     always @(posedge clk) begin
         op_in_2_75 <= op_out_2_74;
         pivot_in_2_75 <= pivot_out_2_74;
         start_in_2_75 <= start_out_2_74;
         swap_in_2_75 <= swap_out_2_74;
     end

     always @(posedge clk) begin
         data_in_2_75 <= data_out_1_75;
     end
  
     processor_AB AB_2_75 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_75),
       .start_in   (start_in_2_75),
       .swap_in   (swap_in_2_75),
       .op_in      (op_in_2_75),
       .pivot_in   (pivot_in_2_75),
       .start_out  (start_out_2_75),
       .swap_out   (swap_out_2_75),
       .data_out   (data_out_2_75),
       .op_out     (op_out_2_75),
       .pivot_out  (pivot_out_2_75),
       .r          (r_2_75)
     );

  // row 2, col 76

     reg start_in_2_76;
     wire start_out_2_76;

     reg swap_in_2_76;
     wire swap_out_2_76;

     reg [1:0] op_in_2_76;
     wire [1:0] op_out_2_76;

     wire r_2_76;

     reg data_in_2_76;
     wire data_out_2_76;

     reg pivot_in_2_76;
     wire pivot_out_2_76;

     always @(posedge clk) begin
         op_in_2_76 <= op_out_2_75;
         pivot_in_2_76 <= pivot_out_2_75;
         start_in_2_76 <= start_out_2_75;
         swap_in_2_76 <= swap_out_2_75;
     end

     always @(posedge clk) begin
         data_in_2_76 <= data_out_1_76;
     end
  
     processor_AB AB_2_76 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_76),
       .start_in   (start_in_2_76),
       .swap_in   (swap_in_2_76),
       .op_in      (op_in_2_76),
       .pivot_in   (pivot_in_2_76),
       .start_out  (start_out_2_76),
       .swap_out   (swap_out_2_76),
       .data_out   (data_out_2_76),
       .op_out     (op_out_2_76),
       .pivot_out  (pivot_out_2_76),
       .r          (r_2_76)
     );

  // row 2, col 77

     reg start_in_2_77;
     wire start_out_2_77;

     reg swap_in_2_77;
     wire swap_out_2_77;

     reg [1:0] op_in_2_77;
     wire [1:0] op_out_2_77;

     wire r_2_77;

     reg data_in_2_77;
     wire data_out_2_77;

     reg pivot_in_2_77;
     wire pivot_out_2_77;

     always @(posedge clk) begin
         op_in_2_77 <= op_out_2_76;
         pivot_in_2_77 <= pivot_out_2_76;
         start_in_2_77 <= start_out_2_76;
         swap_in_2_77 <= swap_out_2_76;
     end

     always @(posedge clk) begin
         data_in_2_77 <= data_out_1_77;
     end
  
     processor_AB AB_2_77 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_77),
       .start_in   (start_in_2_77),
       .swap_in   (swap_in_2_77),
       .op_in      (op_in_2_77),
       .pivot_in   (pivot_in_2_77),
       .start_out  (start_out_2_77),
       .swap_out   (swap_out_2_77),
       .data_out   (data_out_2_77),
       .op_out     (op_out_2_77),
       .pivot_out  (pivot_out_2_77),
       .r          (r_2_77)
     );

  // row 2, col 78

     reg start_in_2_78;
     wire start_out_2_78;

     reg swap_in_2_78;
     wire swap_out_2_78;

     reg [1:0] op_in_2_78;
     wire [1:0] op_out_2_78;

     wire r_2_78;

     reg data_in_2_78;
     wire data_out_2_78;

     reg pivot_in_2_78;
     wire pivot_out_2_78;

     always @(posedge clk) begin
         op_in_2_78 <= op_out_2_77;
         pivot_in_2_78 <= pivot_out_2_77;
         start_in_2_78 <= start_out_2_77;
         swap_in_2_78 <= swap_out_2_77;
     end

     always @(posedge clk) begin
         data_in_2_78 <= data_out_1_78;
     end
  
     processor_AB AB_2_78 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_78),
       .start_in   (start_in_2_78),
       .swap_in   (swap_in_2_78),
       .op_in      (op_in_2_78),
       .pivot_in   (pivot_in_2_78),
       .start_out  (start_out_2_78),
       .swap_out   (swap_out_2_78),
       .data_out   (data_out_2_78),
       .op_out     (op_out_2_78),
       .pivot_out  (pivot_out_2_78),
       .r          (r_2_78)
     );

  // row 2, col 79

     reg start_in_2_79;
     wire start_out_2_79;

     reg swap_in_2_79;
     wire swap_out_2_79;

     reg [1:0] op_in_2_79;
     wire [1:0] op_out_2_79;

     wire r_2_79;

     reg data_in_2_79;
     wire data_out_2_79;

     reg pivot_in_2_79;
     wire pivot_out_2_79;

     always @(posedge clk) begin
         op_in_2_79 <= op_out_2_78;
         pivot_in_2_79 <= pivot_out_2_78;
         start_in_2_79 <= start_out_2_78;
         swap_in_2_79 <= swap_out_2_78;
     end

     always @(posedge clk) begin
         data_in_2_79 <= data_out_1_79;
     end
  
     processor_AB AB_2_79 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_79),
       .start_in   (start_in_2_79),
       .swap_in   (swap_in_2_79),
       .op_in      (op_in_2_79),
       .pivot_in   (pivot_in_2_79),
       .start_out  (start_out_2_79),
       .swap_out   (swap_out_2_79),
       .data_out   (data_out_2_79),
       .op_out     (op_out_2_79),
       .pivot_out  (pivot_out_2_79),
       .r          (r_2_79)
     );

  // row 2, col 80

     reg start_in_2_80;
     wire start_out_2_80;

     reg swap_in_2_80;
     wire swap_out_2_80;

     reg [1:0] op_in_2_80;
     wire [1:0] op_out_2_80;

     wire r_2_80;

     reg data_in_2_80;
     wire data_out_2_80;

     reg pivot_in_2_80;
     wire pivot_out_2_80;

     always @(posedge clk) begin
         op_in_2_80 <= op_out_2_79;
         pivot_in_2_80 <= pivot_out_2_79;
         start_in_2_80 <= start_out_2_79;
         swap_in_2_80 <= swap_out_2_79;
     end

     always @(posedge clk) begin
         data_in_2_80 <= data_out_1_80;
     end
  
     processor_AB AB_2_80 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_80),
       .start_in   (start_in_2_80),
       .swap_in   (swap_in_2_80),
       .op_in      (op_in_2_80),
       .pivot_in   (pivot_in_2_80),
       .start_out  (start_out_2_80),
       .swap_out   (swap_out_2_80),
       .data_out   (data_out_2_80),
       .op_out     (op_out_2_80),
       .pivot_out  (pivot_out_2_80),
       .r          (r_2_80)
     );

  // row 2, col 81

     reg start_in_2_81;
     wire start_out_2_81;

     reg swap_in_2_81;
     wire swap_out_2_81;

     reg [1:0] op_in_2_81;
     wire [1:0] op_out_2_81;

     wire r_2_81;

     reg data_in_2_81;
     wire data_out_2_81;

     reg pivot_in_2_81;
     wire pivot_out_2_81;

     always @(posedge clk) begin
         op_in_2_81 <= op_out_2_80;
         pivot_in_2_81 <= pivot_out_2_80;
         start_in_2_81 <= start_out_2_80;
         swap_in_2_81 <= swap_out_2_80;
     end

     always @(posedge clk) begin
         data_in_2_81 <= data_out_1_81;
     end
  
     processor_AB AB_2_81 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_81),
       .start_in   (start_in_2_81),
       .swap_in   (swap_in_2_81),
       .op_in      (op_in_2_81),
       .pivot_in   (pivot_in_2_81),
       .start_out  (start_out_2_81),
       .swap_out   (swap_out_2_81),
       .data_out   (data_out_2_81),
       .op_out     (op_out_2_81),
       .pivot_out  (pivot_out_2_81),
       .r          (r_2_81)
     );

  // row 2, col 82

     reg start_in_2_82;
     wire start_out_2_82;

     reg swap_in_2_82;
     wire swap_out_2_82;

     reg [1:0] op_in_2_82;
     wire [1:0] op_out_2_82;

     wire r_2_82;

     reg data_in_2_82;
     wire data_out_2_82;

     reg pivot_in_2_82;
     wire pivot_out_2_82;

     always @(posedge clk) begin
         op_in_2_82 <= op_out_2_81;
         pivot_in_2_82 <= pivot_out_2_81;
         start_in_2_82 <= start_out_2_81;
         swap_in_2_82 <= swap_out_2_81;
     end

     always @(posedge clk) begin
         data_in_2_82 <= data_out_1_82;
     end
  
     processor_AB AB_2_82 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_82),
       .start_in   (start_in_2_82),
       .swap_in   (swap_in_2_82),
       .op_in      (op_in_2_82),
       .pivot_in   (pivot_in_2_82),
       .start_out  (start_out_2_82),
       .swap_out   (swap_out_2_82),
       .data_out   (data_out_2_82),
       .op_out     (op_out_2_82),
       .pivot_out  (pivot_out_2_82),
       .r          (r_2_82)
     );

  // row 2, col 83

     reg start_in_2_83;
     wire start_out_2_83;

     reg swap_in_2_83;
     wire swap_out_2_83;

     reg [1:0] op_in_2_83;
     wire [1:0] op_out_2_83;

     wire r_2_83;

     reg data_in_2_83;
     wire data_out_2_83;

     reg pivot_in_2_83;
     wire pivot_out_2_83;

     always @(posedge clk) begin
         op_in_2_83 <= op_out_2_82;
         pivot_in_2_83 <= pivot_out_2_82;
         start_in_2_83 <= start_out_2_82;
         swap_in_2_83 <= swap_out_2_82;
     end

     always @(posedge clk) begin
         data_in_2_83 <= data_out_1_83;
     end
  
     processor_AB AB_2_83 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_83),
       .start_in   (start_in_2_83),
       .swap_in   (swap_in_2_83),
       .op_in      (op_in_2_83),
       .pivot_in   (pivot_in_2_83),
       .start_out  (start_out_2_83),
       .swap_out   (swap_out_2_83),
       .data_out   (data_out_2_83),
       .op_out     (op_out_2_83),
       .pivot_out  (pivot_out_2_83),
       .r          (r_2_83)
     );

  // row 2, col 84

     reg start_in_2_84;
     wire start_out_2_84;

     reg swap_in_2_84;
     wire swap_out_2_84;

     reg [1:0] op_in_2_84;
     wire [1:0] op_out_2_84;

     wire r_2_84;

     reg data_in_2_84;
     wire data_out_2_84;

     reg pivot_in_2_84;
     wire pivot_out_2_84;

     always @(posedge clk) begin
         op_in_2_84 <= op_out_2_83;
         pivot_in_2_84 <= pivot_out_2_83;
         start_in_2_84 <= start_out_2_83;
         swap_in_2_84 <= swap_out_2_83;
     end

     always @(posedge clk) begin
         data_in_2_84 <= data_out_1_84;
     end
  
     processor_AB AB_2_84 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_84),
       .start_in   (start_in_2_84),
       .swap_in   (swap_in_2_84),
       .op_in      (op_in_2_84),
       .pivot_in   (pivot_in_2_84),
       .start_out  (start_out_2_84),
       .swap_out   (swap_out_2_84),
       .data_out   (data_out_2_84),
       .op_out     (op_out_2_84),
       .pivot_out  (pivot_out_2_84),
       .r          (r_2_84)
     );

  // row 2, col 85

     reg start_in_2_85;
     wire start_out_2_85;

     reg swap_in_2_85;
     wire swap_out_2_85;

     reg [1:0] op_in_2_85;
     wire [1:0] op_out_2_85;

     wire r_2_85;

     reg data_in_2_85;
     wire data_out_2_85;

     reg pivot_in_2_85;
     wire pivot_out_2_85;

     always @(posedge clk) begin
         op_in_2_85 <= op_out_2_84;
         pivot_in_2_85 <= pivot_out_2_84;
         start_in_2_85 <= start_out_2_84;
         swap_in_2_85 <= swap_out_2_84;
     end

     always @(posedge clk) begin
         data_in_2_85 <= data_out_1_85;
     end
  
     processor_AB AB_2_85 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_85),
       .start_in   (start_in_2_85),
       .swap_in   (swap_in_2_85),
       .op_in      (op_in_2_85),
       .pivot_in   (pivot_in_2_85),
       .start_out  (start_out_2_85),
       .swap_out   (swap_out_2_85),
       .data_out   (data_out_2_85),
       .op_out     (op_out_2_85),
       .pivot_out  (pivot_out_2_85),
       .r          (r_2_85)
     );

  // row 2, col 86

     reg start_in_2_86;
     wire start_out_2_86;

     reg swap_in_2_86;
     wire swap_out_2_86;

     reg [1:0] op_in_2_86;
     wire [1:0] op_out_2_86;

     wire r_2_86;

     reg data_in_2_86;
     wire data_out_2_86;

     reg pivot_in_2_86;
     wire pivot_out_2_86;

     always @(posedge clk) begin
         op_in_2_86 <= op_out_2_85;
         pivot_in_2_86 <= pivot_out_2_85;
         start_in_2_86 <= start_out_2_85;
         swap_in_2_86 <= swap_out_2_85;
     end

     always @(posedge clk) begin
         data_in_2_86 <= data_out_1_86;
     end
  
     processor_AB AB_2_86 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_86),
       .start_in   (start_in_2_86),
       .swap_in   (swap_in_2_86),
       .op_in      (op_in_2_86),
       .pivot_in   (pivot_in_2_86),
       .start_out  (start_out_2_86),
       .swap_out   (swap_out_2_86),
       .data_out   (data_out_2_86),
       .op_out     (op_out_2_86),
       .pivot_out  (pivot_out_2_86),
       .r          (r_2_86)
     );

  // row 2, col 87

     reg start_in_2_87;
     wire start_out_2_87;

     reg swap_in_2_87;
     wire swap_out_2_87;

     reg [1:0] op_in_2_87;
     wire [1:0] op_out_2_87;

     wire r_2_87;

     reg data_in_2_87;
     wire data_out_2_87;

     reg pivot_in_2_87;
     wire pivot_out_2_87;

     always @(posedge clk) begin
         op_in_2_87 <= op_out_2_86;
         pivot_in_2_87 <= pivot_out_2_86;
         start_in_2_87 <= start_out_2_86;
         swap_in_2_87 <= swap_out_2_86;
     end

     always @(posedge clk) begin
         data_in_2_87 <= data_out_1_87;
     end
  
     processor_AB AB_2_87 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_87),
       .start_in   (start_in_2_87),
       .swap_in   (swap_in_2_87),
       .op_in      (op_in_2_87),
       .pivot_in   (pivot_in_2_87),
       .start_out  (start_out_2_87),
       .swap_out   (swap_out_2_87),
       .data_out   (data_out_2_87),
       .op_out     (op_out_2_87),
       .pivot_out  (pivot_out_2_87),
       .r          (r_2_87)
     );

  // row 2, col 88

     reg start_in_2_88;
     wire start_out_2_88;

     reg swap_in_2_88;
     wire swap_out_2_88;

     reg [1:0] op_in_2_88;
     wire [1:0] op_out_2_88;

     wire r_2_88;

     reg data_in_2_88;
     wire data_out_2_88;

     reg pivot_in_2_88;
     wire pivot_out_2_88;

     always @(posedge clk) begin
         op_in_2_88 <= op_out_2_87;
         pivot_in_2_88 <= pivot_out_2_87;
         start_in_2_88 <= start_out_2_87;
         swap_in_2_88 <= swap_out_2_87;
     end

     always @(posedge clk) begin
         data_in_2_88 <= data_out_1_88;
     end
  
     processor_AB AB_2_88 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_88),
       .start_in   (start_in_2_88),
       .swap_in   (swap_in_2_88),
       .op_in      (op_in_2_88),
       .pivot_in   (pivot_in_2_88),
       .start_out  (start_out_2_88),
       .swap_out   (swap_out_2_88),
       .data_out   (data_out_2_88),
       .op_out     (op_out_2_88),
       .pivot_out  (pivot_out_2_88),
       .r          (r_2_88)
     );

  // row 2, col 89

     reg start_in_2_89;
     wire start_out_2_89;

     reg swap_in_2_89;
     wire swap_out_2_89;

     reg [1:0] op_in_2_89;
     wire [1:0] op_out_2_89;

     wire r_2_89;

     reg data_in_2_89;
     wire data_out_2_89;

     reg pivot_in_2_89;
     wire pivot_out_2_89;

     always @(posedge clk) begin
         op_in_2_89 <= op_out_2_88;
         pivot_in_2_89 <= pivot_out_2_88;
         start_in_2_89 <= start_out_2_88;
         swap_in_2_89 <= swap_out_2_88;
     end

     always @(posedge clk) begin
         data_in_2_89 <= data_out_1_89;
     end
  
     processor_AB AB_2_89 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_89),
       .start_in   (start_in_2_89),
       .swap_in   (swap_in_2_89),
       .op_in      (op_in_2_89),
       .pivot_in   (pivot_in_2_89),
       .start_out  (start_out_2_89),
       .swap_out   (swap_out_2_89),
       .data_out   (data_out_2_89),
       .op_out     (op_out_2_89),
       .pivot_out  (pivot_out_2_89),
       .r          (r_2_89)
     );

  // row 2, col 90

     reg start_in_2_90;
     wire start_out_2_90;

     reg swap_in_2_90;
     wire swap_out_2_90;

     reg [1:0] op_in_2_90;
     wire [1:0] op_out_2_90;

     wire r_2_90;

     reg data_in_2_90;
     wire data_out_2_90;

     reg pivot_in_2_90;
     wire pivot_out_2_90;

     always @(posedge clk) begin
         op_in_2_90 <= op_out_2_89;
         pivot_in_2_90 <= pivot_out_2_89;
         start_in_2_90 <= start_out_2_89;
         swap_in_2_90 <= swap_out_2_89;
     end

     always @(posedge clk) begin
         data_in_2_90 <= data_out_1_90;
     end
  
     processor_AB AB_2_90 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_90),
       .start_in   (start_in_2_90),
       .swap_in   (swap_in_2_90),
       .op_in      (op_in_2_90),
       .pivot_in   (pivot_in_2_90),
       .start_out  (start_out_2_90),
       .swap_out   (swap_out_2_90),
       .data_out   (data_out_2_90),
       .op_out     (op_out_2_90),
       .pivot_out  (pivot_out_2_90),
       .r          (r_2_90)
     );

  // row 2, col 91

     reg start_in_2_91;
     wire start_out_2_91;

     reg swap_in_2_91;
     wire swap_out_2_91;

     reg [1:0] op_in_2_91;
     wire [1:0] op_out_2_91;

     wire r_2_91;

     reg data_in_2_91;
     wire data_out_2_91;

     reg pivot_in_2_91;
     wire pivot_out_2_91;

     always @(posedge clk) begin
         op_in_2_91 <= op_out_2_90;
         pivot_in_2_91 <= pivot_out_2_90;
         start_in_2_91 <= start_out_2_90;
         swap_in_2_91 <= swap_out_2_90;
     end

     always @(posedge clk) begin
         data_in_2_91 <= data_out_1_91;
     end
  
     processor_AB AB_2_91 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_91),
       .start_in   (start_in_2_91),
       .swap_in   (swap_in_2_91),
       .op_in      (op_in_2_91),
       .pivot_in   (pivot_in_2_91),
       .start_out  (start_out_2_91),
       .swap_out   (swap_out_2_91),
       .data_out   (data_out_2_91),
       .op_out     (op_out_2_91),
       .pivot_out  (pivot_out_2_91),
       .r          (r_2_91)
     );

  // row 2, col 92

     reg start_in_2_92;
     wire start_out_2_92;

     reg swap_in_2_92;
     wire swap_out_2_92;

     reg [1:0] op_in_2_92;
     wire [1:0] op_out_2_92;

     wire r_2_92;

     reg data_in_2_92;
     wire data_out_2_92;

     reg pivot_in_2_92;
     wire pivot_out_2_92;

     always @(posedge clk) begin
         op_in_2_92 <= op_out_2_91;
         pivot_in_2_92 <= pivot_out_2_91;
         start_in_2_92 <= start_out_2_91;
         swap_in_2_92 <= swap_out_2_91;
     end

     always @(posedge clk) begin
         data_in_2_92 <= data_out_1_92;
     end
  
     processor_AB AB_2_92 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_92),
       .start_in   (start_in_2_92),
       .swap_in   (swap_in_2_92),
       .op_in      (op_in_2_92),
       .pivot_in   (pivot_in_2_92),
       .start_out  (start_out_2_92),
       .swap_out   (swap_out_2_92),
       .data_out   (data_out_2_92),
       .op_out     (op_out_2_92),
       .pivot_out  (pivot_out_2_92),
       .r          (r_2_92)
     );

  // row 2, col 93

     reg start_in_2_93;
     wire start_out_2_93;

     reg swap_in_2_93;
     wire swap_out_2_93;

     reg [1:0] op_in_2_93;
     wire [1:0] op_out_2_93;

     wire r_2_93;

     reg data_in_2_93;
     wire data_out_2_93;

     reg pivot_in_2_93;
     wire pivot_out_2_93;

     always @(posedge clk) begin
         op_in_2_93 <= op_out_2_92;
         pivot_in_2_93 <= pivot_out_2_92;
         start_in_2_93 <= start_out_2_92;
         swap_in_2_93 <= swap_out_2_92;
     end

     always @(posedge clk) begin
         data_in_2_93 <= data_out_1_93;
     end
  
     processor_AB AB_2_93 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_93),
       .start_in   (start_in_2_93),
       .swap_in   (swap_in_2_93),
       .op_in      (op_in_2_93),
       .pivot_in   (pivot_in_2_93),
       .start_out  (start_out_2_93),
       .swap_out   (swap_out_2_93),
       .data_out   (data_out_2_93),
       .op_out     (op_out_2_93),
       .pivot_out  (pivot_out_2_93),
       .r          (r_2_93)
     );

  // row 2, col 94

     reg start_in_2_94;
     wire start_out_2_94;

     reg swap_in_2_94;
     wire swap_out_2_94;

     reg [1:0] op_in_2_94;
     wire [1:0] op_out_2_94;

     wire r_2_94;

     reg data_in_2_94;
     wire data_out_2_94;

     reg pivot_in_2_94;
     wire pivot_out_2_94;

     always @(posedge clk) begin
         op_in_2_94 <= op_out_2_93;
         pivot_in_2_94 <= pivot_out_2_93;
         start_in_2_94 <= start_out_2_93;
         swap_in_2_94 <= swap_out_2_93;
     end

     always @(posedge clk) begin
         data_in_2_94 <= data_out_1_94;
     end
  
     processor_AB AB_2_94 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_94),
       .start_in   (start_in_2_94),
       .swap_in   (swap_in_2_94),
       .op_in      (op_in_2_94),
       .pivot_in   (pivot_in_2_94),
       .start_out  (start_out_2_94),
       .swap_out   (swap_out_2_94),
       .data_out   (data_out_2_94),
       .op_out     (op_out_2_94),
       .pivot_out  (pivot_out_2_94),
       .r          (r_2_94)
     );

  // row 2, col 95

     reg start_in_2_95;
     wire start_out_2_95;

     reg swap_in_2_95;
     wire swap_out_2_95;

     reg [1:0] op_in_2_95;
     wire [1:0] op_out_2_95;

     wire r_2_95;

     reg data_in_2_95;
     wire data_out_2_95;

     reg pivot_in_2_95;
     wire pivot_out_2_95;

     always @(posedge clk) begin
         op_in_2_95 <= op_out_2_94;
         pivot_in_2_95 <= pivot_out_2_94;
         start_in_2_95 <= start_out_2_94;
         swap_in_2_95 <= swap_out_2_94;
     end

     always @(posedge clk) begin
         data_in_2_95 <= data_out_1_95;
     end
  
     processor_AB AB_2_95 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_95),
       .start_in   (start_in_2_95),
       .swap_in   (swap_in_2_95),
       .op_in      (op_in_2_95),
       .pivot_in   (pivot_in_2_95),
       .start_out  (start_out_2_95),
       .swap_out   (swap_out_2_95),
       .data_out   (data_out_2_95),
       .op_out     (op_out_2_95),
       .pivot_out  (pivot_out_2_95),
       .r          (r_2_95)
     );

  // row 2, col 96

     reg start_in_2_96;
     wire start_out_2_96;

     reg swap_in_2_96;
     wire swap_out_2_96;

     reg [1:0] op_in_2_96;
     wire [1:0] op_out_2_96;

     wire r_2_96;

     reg data_in_2_96;
     wire data_out_2_96;

     reg pivot_in_2_96;
     wire pivot_out_2_96;

     always @(posedge clk) begin
         op_in_2_96 <= op_out_2_95;
         pivot_in_2_96 <= pivot_out_2_95;
         start_in_2_96 <= start_out_2_95;
         swap_in_2_96 <= swap_out_2_95;
     end

     always @(posedge clk) begin
         data_in_2_96 <= data_out_1_96;
     end
  
     processor_AB AB_2_96 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_96),
       .start_in   (start_in_2_96),
       .swap_in   (swap_in_2_96),
       .op_in      (op_in_2_96),
       .pivot_in   (pivot_in_2_96),
       .start_out  (start_out_2_96),
       .swap_out   (swap_out_2_96),
       .data_out   (data_out_2_96),
       .op_out     (op_out_2_96),
       .pivot_out  (pivot_out_2_96),
       .r          (r_2_96)
     );

  // row 2, col 97

     reg start_in_2_97;
     wire start_out_2_97;

     reg swap_in_2_97;
     wire swap_out_2_97;

     reg [1:0] op_in_2_97;
     wire [1:0] op_out_2_97;

     wire r_2_97;

     reg data_in_2_97;
     wire data_out_2_97;

     reg pivot_in_2_97;
     wire pivot_out_2_97;

     always @(posedge clk) begin
         op_in_2_97 <= op_out_2_96;
         pivot_in_2_97 <= pivot_out_2_96;
         start_in_2_97 <= start_out_2_96;
         swap_in_2_97 <= swap_out_2_96;
     end

     always @(posedge clk) begin
         data_in_2_97 <= data_out_1_97;
     end
  
     processor_AB AB_2_97 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_97),
       .start_in   (start_in_2_97),
       .swap_in   (swap_in_2_97),
       .op_in      (op_in_2_97),
       .pivot_in   (pivot_in_2_97),
       .start_out  (start_out_2_97),
       .swap_out   (swap_out_2_97),
       .data_out   (data_out_2_97),
       .op_out     (op_out_2_97),
       .pivot_out  (pivot_out_2_97),
       .r          (r_2_97)
     );

  // row 2, col 98

     reg start_in_2_98;
     wire start_out_2_98;

     reg swap_in_2_98;
     wire swap_out_2_98;

     reg [1:0] op_in_2_98;
     wire [1:0] op_out_2_98;

     wire r_2_98;

     reg data_in_2_98;
     wire data_out_2_98;

     reg pivot_in_2_98;
     wire pivot_out_2_98;

     always @(posedge clk) begin
         op_in_2_98 <= op_out_2_97;
         pivot_in_2_98 <= pivot_out_2_97;
         start_in_2_98 <= start_out_2_97;
         swap_in_2_98 <= swap_out_2_97;
     end

     always @(posedge clk) begin
         data_in_2_98 <= data_out_1_98;
     end
  
     processor_AB AB_2_98 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_98),
       .start_in   (start_in_2_98),
       .swap_in   (swap_in_2_98),
       .op_in      (op_in_2_98),
       .pivot_in   (pivot_in_2_98),
       .start_out  (start_out_2_98),
       .swap_out   (swap_out_2_98),
       .data_out   (data_out_2_98),
       .op_out     (op_out_2_98),
       .pivot_out  (pivot_out_2_98),
       .r          (r_2_98)
     );

  // row 2, col 99

     reg start_in_2_99;
     wire start_out_2_99;

     reg swap_in_2_99;
     wire swap_out_2_99;

     reg [1:0] op_in_2_99;
     wire [1:0] op_out_2_99;

     wire r_2_99;

     reg data_in_2_99;
     wire data_out_2_99;

     reg pivot_in_2_99;
     wire pivot_out_2_99;

     always @(posedge clk) begin
         op_in_2_99 <= op_out_2_98;
         pivot_in_2_99 <= pivot_out_2_98;
         start_in_2_99 <= start_out_2_98;
         swap_in_2_99 <= swap_out_2_98;
     end

     always @(posedge clk) begin
         data_in_2_99 <= data_out_1_99;
     end
  
     processor_AB AB_2_99 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_99),
       .start_in   (start_in_2_99),
       .swap_in   (swap_in_2_99),
       .op_in      (op_in_2_99),
       .pivot_in   (pivot_in_2_99),
       .start_out  (start_out_2_99),
       .swap_out   (swap_out_2_99),
       .data_out   (data_out_2_99),
       .op_out     (op_out_2_99),
       .pivot_out  (pivot_out_2_99),
       .r          (r_2_99)
     );

  // row 2, col 100

     reg start_in_2_100;
     wire start_out_2_100;

     reg swap_in_2_100;
     wire swap_out_2_100;

     reg [1:0] op_in_2_100;
     wire [1:0] op_out_2_100;

     wire r_2_100;

     reg data_in_2_100;
     wire data_out_2_100;

     reg pivot_in_2_100;
     wire pivot_out_2_100;

     always @(posedge clk) begin
         op_in_2_100 <= op_out_2_99;
         pivot_in_2_100 <= pivot_out_2_99;
         start_in_2_100 <= start_out_2_99;
         swap_in_2_100 <= swap_out_2_99;
     end

     always @(posedge clk) begin
         data_in_2_100 <= data_out_1_100;
     end
  
     processor_AB AB_2_100 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_100),
       .start_in   (start_in_2_100),
       .swap_in   (swap_in_2_100),
       .op_in      (op_in_2_100),
       .pivot_in   (pivot_in_2_100),
       .start_out  (start_out_2_100),
       .swap_out   (swap_out_2_100),
       .data_out   (data_out_2_100),
       .op_out     (op_out_2_100),
       .pivot_out  (pivot_out_2_100),
       .r          (r_2_100)
     );

  // row 2, col 101

     reg start_in_2_101;
     wire start_out_2_101;

     reg swap_in_2_101;
     wire swap_out_2_101;

     reg [1:0] op_in_2_101;
     wire [1:0] op_out_2_101;

     wire r_2_101;

     reg data_in_2_101;
     wire data_out_2_101;

     reg pivot_in_2_101;
     wire pivot_out_2_101;

     always @(posedge clk) begin
         op_in_2_101 <= op_out_2_100;
         pivot_in_2_101 <= pivot_out_2_100;
         start_in_2_101 <= start_out_2_100;
         swap_in_2_101 <= swap_out_2_100;
     end

     always @(posedge clk) begin
         data_in_2_101 <= data_out_1_101;
     end
  
     processor_AB AB_2_101 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_101),
       .start_in   (start_in_2_101),
       .swap_in   (swap_in_2_101),
       .op_in      (op_in_2_101),
       .pivot_in   (pivot_in_2_101),
       .start_out  (start_out_2_101),
       .swap_out   (swap_out_2_101),
       .data_out   (data_out_2_101),
       .op_out     (op_out_2_101),
       .pivot_out  (pivot_out_2_101),
       .r          (r_2_101)
     );

  // row 2, col 102

     reg start_in_2_102;
     wire start_out_2_102;

     reg swap_in_2_102;
     wire swap_out_2_102;

     reg [1:0] op_in_2_102;
     wire [1:0] op_out_2_102;

     wire r_2_102;

     reg data_in_2_102;
     wire data_out_2_102;

     reg pivot_in_2_102;
     wire pivot_out_2_102;

     always @(posedge clk) begin
         op_in_2_102 <= op_out_2_101;
         pivot_in_2_102 <= pivot_out_2_101;
         start_in_2_102 <= start_out_2_101;
         swap_in_2_102 <= swap_out_2_101;
     end

     always @(posedge clk) begin
         data_in_2_102 <= data_out_1_102;
     end
  
     processor_AB AB_2_102 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_102),
       .start_in   (start_in_2_102),
       .swap_in   (swap_in_2_102),
       .op_in      (op_in_2_102),
       .pivot_in   (pivot_in_2_102),
       .start_out  (start_out_2_102),
       .swap_out   (swap_out_2_102),
       .data_out   (data_out_2_102),
       .op_out     (op_out_2_102),
       .pivot_out  (pivot_out_2_102),
       .r          (r_2_102)
     );

  // row 2, col 103

     reg start_in_2_103;
     wire start_out_2_103;

     reg swap_in_2_103;
     wire swap_out_2_103;

     reg [1:0] op_in_2_103;
     wire [1:0] op_out_2_103;

     wire r_2_103;

     reg data_in_2_103;
     wire data_out_2_103;

     reg pivot_in_2_103;
     wire pivot_out_2_103;

     always @(posedge clk) begin
         op_in_2_103 <= op_out_2_102;
         pivot_in_2_103 <= pivot_out_2_102;
         start_in_2_103 <= start_out_2_102;
         swap_in_2_103 <= swap_out_2_102;
     end

     always @(posedge clk) begin
         data_in_2_103 <= data_out_1_103;
     end
  
     processor_AB AB_2_103 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_103),
       .start_in   (start_in_2_103),
       .swap_in   (swap_in_2_103),
       .op_in      (op_in_2_103),
       .pivot_in   (pivot_in_2_103),
       .start_out  (start_out_2_103),
       .swap_out   (swap_out_2_103),
       .data_out   (data_out_2_103),
       .op_out     (op_out_2_103),
       .pivot_out  (pivot_out_2_103),
       .r          (r_2_103)
     );

  // row 2, col 104

     reg start_in_2_104;
     wire start_out_2_104;

     reg swap_in_2_104;
     wire swap_out_2_104;

     reg [1:0] op_in_2_104;
     wire [1:0] op_out_2_104;

     wire r_2_104;

     reg data_in_2_104;
     wire data_out_2_104;

     reg pivot_in_2_104;
     wire pivot_out_2_104;

     always @(posedge clk) begin
         op_in_2_104 <= op_out_2_103;
         pivot_in_2_104 <= pivot_out_2_103;
         start_in_2_104 <= start_out_2_103;
         swap_in_2_104 <= swap_out_2_103;
     end

     always @(posedge clk) begin
         data_in_2_104 <= data_out_1_104;
     end
  
     processor_AB AB_2_104 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_104),
       .start_in   (start_in_2_104),
       .swap_in   (swap_in_2_104),
       .op_in      (op_in_2_104),
       .pivot_in   (pivot_in_2_104),
       .start_out  (start_out_2_104),
       .swap_out   (swap_out_2_104),
       .data_out   (data_out_2_104),
       .op_out     (op_out_2_104),
       .pivot_out  (pivot_out_2_104),
       .r          (r_2_104)
     );

  // row 2, col 105

     reg start_in_2_105;
     wire start_out_2_105;

     reg swap_in_2_105;
     wire swap_out_2_105;

     reg [1:0] op_in_2_105;
     wire [1:0] op_out_2_105;

     wire r_2_105;

     reg data_in_2_105;
     wire data_out_2_105;

     reg pivot_in_2_105;
     wire pivot_out_2_105;

     always @(posedge clk) begin
         op_in_2_105 <= op_out_2_104;
         pivot_in_2_105 <= pivot_out_2_104;
         start_in_2_105 <= start_out_2_104;
         swap_in_2_105 <= swap_out_2_104;
     end

     always @(posedge clk) begin
         data_in_2_105 <= data_out_1_105;
     end
  
     processor_AB AB_2_105 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_105),
       .start_in   (start_in_2_105),
       .swap_in   (swap_in_2_105),
       .op_in      (op_in_2_105),
       .pivot_in   (pivot_in_2_105),
       .start_out  (start_out_2_105),
       .swap_out   (swap_out_2_105),
       .data_out   (data_out_2_105),
       .op_out     (op_out_2_105),
       .pivot_out  (pivot_out_2_105),
       .r          (r_2_105)
     );

  // row 2, col 106

     reg start_in_2_106;
     wire start_out_2_106;

     reg swap_in_2_106;
     wire swap_out_2_106;

     reg [1:0] op_in_2_106;
     wire [1:0] op_out_2_106;

     wire r_2_106;

     reg data_in_2_106;
     wire data_out_2_106;

     reg pivot_in_2_106;
     wire pivot_out_2_106;

     always @(posedge clk) begin
         op_in_2_106 <= op_out_2_105;
         pivot_in_2_106 <= pivot_out_2_105;
         start_in_2_106 <= start_out_2_105;
         swap_in_2_106 <= swap_out_2_105;
     end

     always @(posedge clk) begin
         data_in_2_106 <= data_out_1_106;
     end
  
     processor_AB AB_2_106 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_106),
       .start_in   (start_in_2_106),
       .swap_in   (swap_in_2_106),
       .op_in      (op_in_2_106),
       .pivot_in   (pivot_in_2_106),
       .start_out  (start_out_2_106),
       .swap_out   (swap_out_2_106),
       .data_out   (data_out_2_106),
       .op_out     (op_out_2_106),
       .pivot_out  (pivot_out_2_106),
       .r          (r_2_106)
     );

  // row 2, col 107

     reg start_in_2_107;
     wire start_out_2_107;

     reg swap_in_2_107;
     wire swap_out_2_107;

     reg [1:0] op_in_2_107;
     wire [1:0] op_out_2_107;

     wire r_2_107;

     reg data_in_2_107;
     wire data_out_2_107;

     reg pivot_in_2_107;
     wire pivot_out_2_107;

     always @(posedge clk) begin
         op_in_2_107 <= op_out_2_106;
         pivot_in_2_107 <= pivot_out_2_106;
         start_in_2_107 <= start_out_2_106;
         swap_in_2_107 <= swap_out_2_106;
     end

     always @(posedge clk) begin
         data_in_2_107 <= data_out_1_107;
     end
  
     processor_AB AB_2_107 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_107),
       .start_in   (start_in_2_107),
       .swap_in   (swap_in_2_107),
       .op_in      (op_in_2_107),
       .pivot_in   (pivot_in_2_107),
       .start_out  (start_out_2_107),
       .swap_out   (swap_out_2_107),
       .data_out   (data_out_2_107),
       .op_out     (op_out_2_107),
       .pivot_out  (pivot_out_2_107),
       .r          (r_2_107)
     );

  // row 2, col 108

     reg start_in_2_108;
     wire start_out_2_108;

     reg swap_in_2_108;
     wire swap_out_2_108;

     reg [1:0] op_in_2_108;
     wire [1:0] op_out_2_108;

     wire r_2_108;

     reg data_in_2_108;
     wire data_out_2_108;

     reg pivot_in_2_108;
     wire pivot_out_2_108;

     always @(posedge clk) begin
         op_in_2_108 <= op_out_2_107;
         pivot_in_2_108 <= pivot_out_2_107;
         start_in_2_108 <= start_out_2_107;
         swap_in_2_108 <= swap_out_2_107;
     end

     always @(posedge clk) begin
         data_in_2_108 <= data_out_1_108;
     end
  
     processor_AB AB_2_108 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_108),
       .start_in   (start_in_2_108),
       .swap_in   (swap_in_2_108),
       .op_in      (op_in_2_108),
       .pivot_in   (pivot_in_2_108),
       .start_out  (start_out_2_108),
       .swap_out   (swap_out_2_108),
       .data_out   (data_out_2_108),
       .op_out     (op_out_2_108),
       .pivot_out  (pivot_out_2_108),
       .r          (r_2_108)
     );

  // row 2, col 109

     reg start_in_2_109;
     wire start_out_2_109;

     reg swap_in_2_109;
     wire swap_out_2_109;

     reg [1:0] op_in_2_109;
     wire [1:0] op_out_2_109;

     wire r_2_109;

     reg data_in_2_109;
     wire data_out_2_109;

     reg pivot_in_2_109;
     wire pivot_out_2_109;

     always @(posedge clk) begin
         op_in_2_109 <= op_out_2_108;
         pivot_in_2_109 <= pivot_out_2_108;
         start_in_2_109 <= start_out_2_108;
         swap_in_2_109 <= swap_out_2_108;
     end

     always @(posedge clk) begin
         data_in_2_109 <= data_out_1_109;
     end
  
     processor_AB AB_2_109 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_109),
       .start_in   (start_in_2_109),
       .swap_in   (swap_in_2_109),
       .op_in      (op_in_2_109),
       .pivot_in   (pivot_in_2_109),
       .start_out  (start_out_2_109),
       .swap_out   (swap_out_2_109),
       .data_out   (data_out_2_109),
       .op_out     (op_out_2_109),
       .pivot_out  (pivot_out_2_109),
       .r          (r_2_109)
     );

  // row 2, col 110

     reg start_in_2_110;
     wire start_out_2_110;

     reg swap_in_2_110;
     wire swap_out_2_110;

     reg [1:0] op_in_2_110;
     wire [1:0] op_out_2_110;

     wire r_2_110;

     reg data_in_2_110;
     wire data_out_2_110;

     reg pivot_in_2_110;
     wire pivot_out_2_110;

     always @(posedge clk) begin
         op_in_2_110 <= op_out_2_109;
         pivot_in_2_110 <= pivot_out_2_109;
         start_in_2_110 <= start_out_2_109;
         swap_in_2_110 <= swap_out_2_109;
     end

     always @(posedge clk) begin
         data_in_2_110 <= data_out_1_110;
     end
  
     processor_AB AB_2_110 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_110),
       .start_in   (start_in_2_110),
       .swap_in   (swap_in_2_110),
       .op_in      (op_in_2_110),
       .pivot_in   (pivot_in_2_110),
       .start_out  (start_out_2_110),
       .swap_out   (swap_out_2_110),
       .data_out   (data_out_2_110),
       .op_out     (op_out_2_110),
       .pivot_out  (pivot_out_2_110),
       .r          (r_2_110)
     );

  // row 2, col 111

     reg start_in_2_111;
     wire start_out_2_111;

     reg swap_in_2_111;
     wire swap_out_2_111;

     reg [1:0] op_in_2_111;
     wire [1:0] op_out_2_111;

     wire r_2_111;

     reg data_in_2_111;
     wire data_out_2_111;

     reg pivot_in_2_111;
     wire pivot_out_2_111;

     always @(posedge clk) begin
         op_in_2_111 <= op_out_2_110;
         pivot_in_2_111 <= pivot_out_2_110;
         start_in_2_111 <= start_out_2_110;
         swap_in_2_111 <= swap_out_2_110;
     end

     always @(posedge clk) begin
         data_in_2_111 <= data_out_1_111;
     end
  
     processor_AB AB_2_111 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_111),
       .start_in   (start_in_2_111),
       .swap_in   (swap_in_2_111),
       .op_in      (op_in_2_111),
       .pivot_in   (pivot_in_2_111),
       .start_out  (start_out_2_111),
       .swap_out   (swap_out_2_111),
       .data_out   (data_out_2_111),
       .op_out     (op_out_2_111),
       .pivot_out  (pivot_out_2_111),
       .r          (r_2_111)
     );

  // row 2, col 112

     reg start_in_2_112;
     wire start_out_2_112;

     reg swap_in_2_112;
     wire swap_out_2_112;

     reg [1:0] op_in_2_112;
     wire [1:0] op_out_2_112;

     wire r_2_112;

     reg data_in_2_112;
     wire data_out_2_112;

     reg pivot_in_2_112;
     wire pivot_out_2_112;

     always @(posedge clk) begin
         op_in_2_112 <= op_out_2_111;
         pivot_in_2_112 <= pivot_out_2_111;
         start_in_2_112 <= start_out_2_111;
         swap_in_2_112 <= swap_out_2_111;
     end

     always @(posedge clk) begin
         data_in_2_112 <= data_out_1_112;
     end
  
     processor_AB AB_2_112 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_112),
       .start_in   (start_in_2_112),
       .swap_in   (swap_in_2_112),
       .op_in      (op_in_2_112),
       .pivot_in   (pivot_in_2_112),
       .start_out  (start_out_2_112),
       .swap_out   (swap_out_2_112),
       .data_out   (data_out_2_112),
       .op_out     (op_out_2_112),
       .pivot_out  (pivot_out_2_112),
       .r          (r_2_112)
     );

  // row 2, col 113

     reg start_in_2_113;
     wire start_out_2_113;

     reg swap_in_2_113;
     wire swap_out_2_113;

     reg [1:0] op_in_2_113;
     wire [1:0] op_out_2_113;

     wire r_2_113;

     reg data_in_2_113;
     wire data_out_2_113;

     reg pivot_in_2_113;
     wire pivot_out_2_113;

     always @(posedge clk) begin
         op_in_2_113 <= op_out_2_112;
         pivot_in_2_113 <= pivot_out_2_112;
         start_in_2_113 <= start_out_2_112;
         swap_in_2_113 <= swap_out_2_112;
     end

     always @(posedge clk) begin
         data_in_2_113 <= data_out_1_113;
     end
  
     processor_AB AB_2_113 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_113),
       .start_in   (start_in_2_113),
       .swap_in   (swap_in_2_113),
       .op_in      (op_in_2_113),
       .pivot_in   (pivot_in_2_113),
       .start_out  (start_out_2_113),
       .swap_out   (swap_out_2_113),
       .data_out   (data_out_2_113),
       .op_out     (op_out_2_113),
       .pivot_out  (pivot_out_2_113),
       .r          (r_2_113)
     );

  // row 2, col 114

     reg start_in_2_114;
     wire start_out_2_114;

     reg swap_in_2_114;
     wire swap_out_2_114;

     reg [1:0] op_in_2_114;
     wire [1:0] op_out_2_114;

     wire r_2_114;

     reg data_in_2_114;
     wire data_out_2_114;

     reg pivot_in_2_114;
     wire pivot_out_2_114;

     always @(posedge clk) begin
         op_in_2_114 <= op_out_2_113;
         pivot_in_2_114 <= pivot_out_2_113;
         start_in_2_114 <= start_out_2_113;
         swap_in_2_114 <= swap_out_2_113;
     end

     always @(posedge clk) begin
         data_in_2_114 <= data_out_1_114;
     end
  
     processor_AB AB_2_114 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_114),
       .start_in   (start_in_2_114),
       .swap_in   (swap_in_2_114),
       .op_in      (op_in_2_114),
       .pivot_in   (pivot_in_2_114),
       .start_out  (start_out_2_114),
       .swap_out   (swap_out_2_114),
       .data_out   (data_out_2_114),
       .op_out     (op_out_2_114),
       .pivot_out  (pivot_out_2_114),
       .r          (r_2_114)
     );

  // row 2, col 115

     reg start_in_2_115;
     wire start_out_2_115;

     reg swap_in_2_115;
     wire swap_out_2_115;

     reg [1:0] op_in_2_115;
     wire [1:0] op_out_2_115;

     wire r_2_115;

     reg data_in_2_115;
     wire data_out_2_115;

     reg pivot_in_2_115;
     wire pivot_out_2_115;

     always @(posedge clk) begin
         op_in_2_115 <= op_out_2_114;
         pivot_in_2_115 <= pivot_out_2_114;
         start_in_2_115 <= start_out_2_114;
         swap_in_2_115 <= swap_out_2_114;
     end

     always @(posedge clk) begin
         data_in_2_115 <= data_out_1_115;
     end
  
     processor_AB AB_2_115 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_115),
       .start_in   (start_in_2_115),
       .swap_in   (swap_in_2_115),
       .op_in      (op_in_2_115),
       .pivot_in   (pivot_in_2_115),
       .start_out  (start_out_2_115),
       .swap_out   (swap_out_2_115),
       .data_out   (data_out_2_115),
       .op_out     (op_out_2_115),
       .pivot_out  (pivot_out_2_115),
       .r          (r_2_115)
     );

  // row 2, col 116

     reg start_in_2_116;
     wire start_out_2_116;

     reg swap_in_2_116;
     wire swap_out_2_116;

     reg [1:0] op_in_2_116;
     wire [1:0] op_out_2_116;

     wire r_2_116;

     reg data_in_2_116;
     wire data_out_2_116;

     reg pivot_in_2_116;
     wire pivot_out_2_116;

     always @(posedge clk) begin
         op_in_2_116 <= op_out_2_115;
         pivot_in_2_116 <= pivot_out_2_115;
         start_in_2_116 <= start_out_2_115;
         swap_in_2_116 <= swap_out_2_115;
     end

     always @(posedge clk) begin
         data_in_2_116 <= data_out_1_116;
     end
  
     processor_AB AB_2_116 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_116),
       .start_in   (start_in_2_116),
       .swap_in   (swap_in_2_116),
       .op_in      (op_in_2_116),
       .pivot_in   (pivot_in_2_116),
       .start_out  (start_out_2_116),
       .swap_out   (swap_out_2_116),
       .data_out   (data_out_2_116),
       .op_out     (op_out_2_116),
       .pivot_out  (pivot_out_2_116),
       .r          (r_2_116)
     );

  // row 2, col 117

     reg start_in_2_117;
     wire start_out_2_117;

     reg swap_in_2_117;
     wire swap_out_2_117;

     reg [1:0] op_in_2_117;
     wire [1:0] op_out_2_117;

     wire r_2_117;

     reg data_in_2_117;
     wire data_out_2_117;

     reg pivot_in_2_117;
     wire pivot_out_2_117;

     always @(posedge clk) begin
         op_in_2_117 <= op_out_2_116;
         pivot_in_2_117 <= pivot_out_2_116;
         start_in_2_117 <= start_out_2_116;
         swap_in_2_117 <= swap_out_2_116;
     end

     always @(posedge clk) begin
         data_in_2_117 <= data_out_1_117;
     end
  
     processor_AB AB_2_117 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_117),
       .start_in   (start_in_2_117),
       .swap_in   (swap_in_2_117),
       .op_in      (op_in_2_117),
       .pivot_in   (pivot_in_2_117),
       .start_out  (start_out_2_117),
       .swap_out   (swap_out_2_117),
       .data_out   (data_out_2_117),
       .op_out     (op_out_2_117),
       .pivot_out  (pivot_out_2_117),
       .r          (r_2_117)
     );

  // row 2, col 118

     reg start_in_2_118;
     wire start_out_2_118;

     reg swap_in_2_118;
     wire swap_out_2_118;

     reg [1:0] op_in_2_118;
     wire [1:0] op_out_2_118;

     wire r_2_118;

     reg data_in_2_118;
     wire data_out_2_118;

     reg pivot_in_2_118;
     wire pivot_out_2_118;

     always @(posedge clk) begin
         op_in_2_118 <= op_out_2_117;
         pivot_in_2_118 <= pivot_out_2_117;
         start_in_2_118 <= start_out_2_117;
         swap_in_2_118 <= swap_out_2_117;
     end

     always @(posedge clk) begin
         data_in_2_118 <= data_out_1_118;
     end
  
     processor_AB AB_2_118 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_118),
       .start_in   (start_in_2_118),
       .swap_in   (swap_in_2_118),
       .op_in      (op_in_2_118),
       .pivot_in   (pivot_in_2_118),
       .start_out  (start_out_2_118),
       .swap_out   (swap_out_2_118),
       .data_out   (data_out_2_118),
       .op_out     (op_out_2_118),
       .pivot_out  (pivot_out_2_118),
       .r          (r_2_118)
     );

  // row 2, col 119

     reg start_in_2_119;
     wire start_out_2_119;

     reg swap_in_2_119;
     wire swap_out_2_119;

     reg [1:0] op_in_2_119;
     wire [1:0] op_out_2_119;

     wire r_2_119;

     reg data_in_2_119;
     wire data_out_2_119;

     reg pivot_in_2_119;
     wire pivot_out_2_119;

     always @(posedge clk) begin
         op_in_2_119 <= op_out_2_118;
         pivot_in_2_119 <= pivot_out_2_118;
         start_in_2_119 <= start_out_2_118;
         swap_in_2_119 <= swap_out_2_118;
     end

     always @(posedge clk) begin
         data_in_2_119 <= data_out_1_119;
     end
  
     processor_AB AB_2_119 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_119),
       .start_in   (start_in_2_119),
       .swap_in   (swap_in_2_119),
       .op_in      (op_in_2_119),
       .pivot_in   (pivot_in_2_119),
       .start_out  (start_out_2_119),
       .swap_out   (swap_out_2_119),
       .data_out   (data_out_2_119),
       .op_out     (op_out_2_119),
       .pivot_out  (pivot_out_2_119),
       .r          (r_2_119)
     );

  // row 2, col 120

     reg start_in_2_120;
     wire start_out_2_120;

     reg swap_in_2_120;
     wire swap_out_2_120;

     reg [1:0] op_in_2_120;
     wire [1:0] op_out_2_120;

     wire r_2_120;

     reg data_in_2_120;
     wire data_out_2_120;

     reg pivot_in_2_120;
     wire pivot_out_2_120;

     always @(posedge clk) begin
         op_in_2_120 <= op_out_2_119;
         pivot_in_2_120 <= pivot_out_2_119;
         start_in_2_120 <= start_out_2_119;
         swap_in_2_120 <= swap_out_2_119;
     end

     always @(posedge clk) begin
         data_in_2_120 <= data_out_1_120;
     end
  
     processor_AB AB_2_120 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_120),
       .start_in   (start_in_2_120),
       .swap_in   (swap_in_2_120),
       .op_in      (op_in_2_120),
       .pivot_in   (pivot_in_2_120),
       .start_out  (start_out_2_120),
       .swap_out   (swap_out_2_120),
       .data_out   (data_out_2_120),
       .op_out     (op_out_2_120),
       .pivot_out  (pivot_out_2_120),
       .r          (r_2_120)
     );

  // row 2, col 121

     reg start_in_2_121;
     wire start_out_2_121;

     reg swap_in_2_121;
     wire swap_out_2_121;

     reg [1:0] op_in_2_121;
     wire [1:0] op_out_2_121;

     wire r_2_121;

     reg data_in_2_121;
     wire data_out_2_121;

     reg pivot_in_2_121;
     wire pivot_out_2_121;

     always @(posedge clk) begin
         op_in_2_121 <= op_out_2_120;
         pivot_in_2_121 <= pivot_out_2_120;
         start_in_2_121 <= start_out_2_120;
         swap_in_2_121 <= swap_out_2_120;
     end

     always @(posedge clk) begin
         data_in_2_121 <= data_out_1_121;
     end
  
     processor_AB AB_2_121 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_121),
       .start_in   (start_in_2_121),
       .swap_in   (swap_in_2_121),
       .op_in      (op_in_2_121),
       .pivot_in   (pivot_in_2_121),
       .start_out  (start_out_2_121),
       .swap_out   (swap_out_2_121),
       .data_out   (data_out_2_121),
       .op_out     (op_out_2_121),
       .pivot_out  (pivot_out_2_121),
       .r          (r_2_121)
     );

  // row 2, col 122

     reg start_in_2_122;
     wire start_out_2_122;

     reg swap_in_2_122;
     wire swap_out_2_122;

     reg [1:0] op_in_2_122;
     wire [1:0] op_out_2_122;

     wire r_2_122;

     reg data_in_2_122;
     wire data_out_2_122;

     reg pivot_in_2_122;
     wire pivot_out_2_122;

     always @(posedge clk) begin
         op_in_2_122 <= op_out_2_121;
         pivot_in_2_122 <= pivot_out_2_121;
         start_in_2_122 <= start_out_2_121;
         swap_in_2_122 <= swap_out_2_121;
     end

     always @(posedge clk) begin
         data_in_2_122 <= data_out_1_122;
     end
  
     processor_AB AB_2_122 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_122),
       .start_in   (start_in_2_122),
       .swap_in   (swap_in_2_122),
       .op_in      (op_in_2_122),
       .pivot_in   (pivot_in_2_122),
       .start_out  (start_out_2_122),
       .swap_out   (swap_out_2_122),
       .data_out   (data_out_2_122),
       .op_out     (op_out_2_122),
       .pivot_out  (pivot_out_2_122),
       .r          (r_2_122)
     );

  // row 2, col 123

     reg start_in_2_123;
     wire start_out_2_123;

     reg swap_in_2_123;
     wire swap_out_2_123;

     reg [1:0] op_in_2_123;
     wire [1:0] op_out_2_123;

     wire r_2_123;

     reg data_in_2_123;
     wire data_out_2_123;

     reg pivot_in_2_123;
     wire pivot_out_2_123;

     always @(posedge clk) begin
         op_in_2_123 <= op_out_2_122;
         pivot_in_2_123 <= pivot_out_2_122;
         start_in_2_123 <= start_out_2_122;
         swap_in_2_123 <= swap_out_2_122;
     end

     always @(posedge clk) begin
         data_in_2_123 <= data_out_1_123;
     end
  
     processor_AB AB_2_123 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_123),
       .start_in   (start_in_2_123),
       .swap_in   (swap_in_2_123),
       .op_in      (op_in_2_123),
       .pivot_in   (pivot_in_2_123),
       .start_out  (start_out_2_123),
       .swap_out   (swap_out_2_123),
       .data_out   (data_out_2_123),
       .op_out     (op_out_2_123),
       .pivot_out  (pivot_out_2_123),
       .r          (r_2_123)
     );

  // row 2, col 124

     reg start_in_2_124;
     wire start_out_2_124;

     reg swap_in_2_124;
     wire swap_out_2_124;

     reg [1:0] op_in_2_124;
     wire [1:0] op_out_2_124;

     wire r_2_124;

     reg data_in_2_124;
     wire data_out_2_124;

     reg pivot_in_2_124;
     wire pivot_out_2_124;

     always @(posedge clk) begin
         op_in_2_124 <= op_out_2_123;
         pivot_in_2_124 <= pivot_out_2_123;
         start_in_2_124 <= start_out_2_123;
         swap_in_2_124 <= swap_out_2_123;
     end

     always @(posedge clk) begin
         data_in_2_124 <= data_out_1_124;
     end
  
     processor_AB AB_2_124 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_124),
       .start_in   (start_in_2_124),
       .swap_in   (swap_in_2_124),
       .op_in      (op_in_2_124),
       .pivot_in   (pivot_in_2_124),
       .start_out  (start_out_2_124),
       .swap_out   (swap_out_2_124),
       .data_out   (data_out_2_124),
       .op_out     (op_out_2_124),
       .pivot_out  (pivot_out_2_124),
       .r          (r_2_124)
     );

  // row 2, col 125

     reg start_in_2_125;
     wire start_out_2_125;

     reg swap_in_2_125;
     wire swap_out_2_125;

     reg [1:0] op_in_2_125;
     wire [1:0] op_out_2_125;

     wire r_2_125;

     reg data_in_2_125;
     wire data_out_2_125;

     reg pivot_in_2_125;
     wire pivot_out_2_125;

     always @(posedge clk) begin
         op_in_2_125 <= op_out_2_124;
         pivot_in_2_125 <= pivot_out_2_124;
         start_in_2_125 <= start_out_2_124;
         swap_in_2_125 <= swap_out_2_124;
     end

     always @(posedge clk) begin
         data_in_2_125 <= data_out_1_125;
     end
  
     processor_AB AB_2_125 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_125),
       .start_in   (start_in_2_125),
       .swap_in   (swap_in_2_125),
       .op_in      (op_in_2_125),
       .pivot_in   (pivot_in_2_125),
       .start_out  (start_out_2_125),
       .swap_out   (swap_out_2_125),
       .data_out   (data_out_2_125),
       .op_out     (op_out_2_125),
       .pivot_out  (pivot_out_2_125),
       .r          (r_2_125)
     );

  // row 2, col 126

     reg start_in_2_126;
     wire start_out_2_126;

     reg swap_in_2_126;
     wire swap_out_2_126;

     reg [1:0] op_in_2_126;
     wire [1:0] op_out_2_126;

     wire r_2_126;

     reg data_in_2_126;
     wire data_out_2_126;

     reg pivot_in_2_126;
     wire pivot_out_2_126;

     always @(posedge clk) begin
         op_in_2_126 <= op_out_2_125;
         pivot_in_2_126 <= pivot_out_2_125;
         start_in_2_126 <= start_out_2_125;
         swap_in_2_126 <= swap_out_2_125;
     end

     always @(posedge clk) begin
         data_in_2_126 <= data_out_1_126;
     end
  
     processor_AB AB_2_126 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_126),
       .start_in   (start_in_2_126),
       .swap_in   (swap_in_2_126),
       .op_in      (op_in_2_126),
       .pivot_in   (pivot_in_2_126),
       .start_out  (start_out_2_126),
       .swap_out   (swap_out_2_126),
       .data_out   (data_out_2_126),
       .op_out     (op_out_2_126),
       .pivot_out  (pivot_out_2_126),
       .r          (r_2_126)
     );

  // row 2, col 127

     reg start_in_2_127;
     wire start_out_2_127;

     reg swap_in_2_127;
     wire swap_out_2_127;

     reg [1:0] op_in_2_127;
     wire [1:0] op_out_2_127;

     wire r_2_127;

     reg data_in_2_127;
     wire data_out_2_127;

     reg pivot_in_2_127;
     wire pivot_out_2_127;

     always @(posedge clk) begin
         op_in_2_127 <= op_out_2_126;
         pivot_in_2_127 <= pivot_out_2_126;
         start_in_2_127 <= start_out_2_126;
         swap_in_2_127 <= swap_out_2_126;
     end

     always @(posedge clk) begin
         data_in_2_127 <= data_out_1_127;
     end
  
     processor_AB AB_2_127 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_127),
       .start_in   (start_in_2_127),
       .swap_in   (swap_in_2_127),
       .op_in      (op_in_2_127),
       .pivot_in   (pivot_in_2_127),
       .start_out  (start_out_2_127),
       .swap_out   (swap_out_2_127),
       .data_out   (data_out_2_127),
       .op_out     (op_out_2_127),
       .pivot_out  (pivot_out_2_127),
       .r          (r_2_127)
     );

  // row 2, col 128

     reg start_in_2_128;
     wire start_out_2_128;

     reg swap_in_2_128;
     wire swap_out_2_128;

     reg [1:0] op_in_2_128;
     wire [1:0] op_out_2_128;

     wire r_2_128;

     reg data_in_2_128;
     wire data_out_2_128;

     reg pivot_in_2_128;
     wire pivot_out_2_128;

     always @(posedge clk) begin
         op_in_2_128 <= op_out_2_127;
         pivot_in_2_128 <= pivot_out_2_127;
         start_in_2_128 <= start_out_2_127;
         swap_in_2_128 <= swap_out_2_127;
     end

     always @(posedge clk) begin
         data_in_2_128 <= data_out_1_128;
     end
  
     processor_AB AB_2_128 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_128),
       .start_in   (start_in_2_128),
       .swap_in   (swap_in_2_128),
       .op_in      (op_in_2_128),
       .pivot_in   (pivot_in_2_128),
       .start_out  (start_out_2_128),
       .swap_out   (swap_out_2_128),
       .data_out   (data_out_2_128),
       .op_out     (op_out_2_128),
       .pivot_out  (pivot_out_2_128),
       .r          (r_2_128)
     );

  // row 2, col 129

     reg start_in_2_129;
     wire start_out_2_129;

     reg swap_in_2_129;
     wire swap_out_2_129;

     reg [1:0] op_in_2_129;
     wire [1:0] op_out_2_129;

     wire r_2_129;

     reg data_in_2_129;
     wire data_out_2_129;

     reg pivot_in_2_129;
     wire pivot_out_2_129;

     always @(posedge clk) begin
         op_in_2_129 <= op_out_2_128;
         pivot_in_2_129 <= pivot_out_2_128;
         start_in_2_129 <= start_out_2_128;
         swap_in_2_129 <= swap_out_2_128;
     end

     always @(posedge clk) begin
         data_in_2_129 <= data_out_1_129;
     end
  
     processor_AB AB_2_129 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_129),
       .start_in   (start_in_2_129),
       .swap_in   (swap_in_2_129),
       .op_in      (op_in_2_129),
       .pivot_in   (pivot_in_2_129),
       .start_out  (start_out_2_129),
       .swap_out   (swap_out_2_129),
       .data_out   (data_out_2_129),
       .op_out     (op_out_2_129),
       .pivot_out  (pivot_out_2_129),
       .r          (r_2_129)
     );

  // row 2, col 130

     reg start_in_2_130;
     wire start_out_2_130;

     reg swap_in_2_130;
     wire swap_out_2_130;

     reg [1:0] op_in_2_130;
     wire [1:0] op_out_2_130;

     wire r_2_130;

     reg data_in_2_130;
     wire data_out_2_130;

     reg pivot_in_2_130;
     wire pivot_out_2_130;

     always @(posedge clk) begin
         op_in_2_130 <= op_out_2_129;
         pivot_in_2_130 <= pivot_out_2_129;
         start_in_2_130 <= start_out_2_129;
         swap_in_2_130 <= swap_out_2_129;
     end

     always @(posedge clk) begin
         data_in_2_130 <= data_out_1_130;
     end
  
     processor_AB AB_2_130 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_130),
       .start_in   (start_in_2_130),
       .swap_in   (swap_in_2_130),
       .op_in      (op_in_2_130),
       .pivot_in   (pivot_in_2_130),
       .start_out  (start_out_2_130),
       .swap_out   (swap_out_2_130),
       .data_out   (data_out_2_130),
       .op_out     (op_out_2_130),
       .pivot_out  (pivot_out_2_130),
       .r          (r_2_130)
     );

  // row 2, col 131

     reg start_in_2_131;
     wire start_out_2_131;

     reg swap_in_2_131;
     wire swap_out_2_131;

     reg [1:0] op_in_2_131;
     wire [1:0] op_out_2_131;

     wire r_2_131;

     reg data_in_2_131;
     wire data_out_2_131;

     reg pivot_in_2_131;
     wire pivot_out_2_131;

     always @(posedge clk) begin
         op_in_2_131 <= op_out_2_130;
         pivot_in_2_131 <= pivot_out_2_130;
         start_in_2_131 <= start_out_2_130;
         swap_in_2_131 <= swap_out_2_130;
     end

     always @(posedge clk) begin
         data_in_2_131 <= data_out_1_131;
     end
  
     processor_AB AB_2_131 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_131),
       .start_in   (start_in_2_131),
       .swap_in   (swap_in_2_131),
       .op_in      (op_in_2_131),
       .pivot_in   (pivot_in_2_131),
       .start_out  (start_out_2_131),
       .swap_out   (swap_out_2_131),
       .data_out   (data_out_2_131),
       .op_out     (op_out_2_131),
       .pivot_out  (pivot_out_2_131),
       .r          (r_2_131)
     );

  // row 2, col 132

     reg start_in_2_132;
     wire start_out_2_132;

     reg swap_in_2_132;
     wire swap_out_2_132;

     reg [1:0] op_in_2_132;
     wire [1:0] op_out_2_132;

     wire r_2_132;

     reg data_in_2_132;
     wire data_out_2_132;

     reg pivot_in_2_132;
     wire pivot_out_2_132;

     always @(posedge clk) begin
         op_in_2_132 <= op_out_2_131;
         pivot_in_2_132 <= pivot_out_2_131;
         start_in_2_132 <= start_out_2_131;
         swap_in_2_132 <= swap_out_2_131;
     end

     always @(posedge clk) begin
         data_in_2_132 <= data_out_1_132;
     end
  
     processor_AB AB_2_132 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_132),
       .start_in   (start_in_2_132),
       .swap_in   (swap_in_2_132),
       .op_in      (op_in_2_132),
       .pivot_in   (pivot_in_2_132),
       .start_out  (start_out_2_132),
       .swap_out   (swap_out_2_132),
       .data_out   (data_out_2_132),
       .op_out     (op_out_2_132),
       .pivot_out  (pivot_out_2_132),
       .r          (r_2_132)
     );

  // row 2, col 133

     reg start_in_2_133;
     wire start_out_2_133;

     reg swap_in_2_133;
     wire swap_out_2_133;

     reg [1:0] op_in_2_133;
     wire [1:0] op_out_2_133;

     wire r_2_133;

     reg data_in_2_133;
     wire data_out_2_133;

     reg pivot_in_2_133;
     wire pivot_out_2_133;

     always @(posedge clk) begin
         op_in_2_133 <= op_out_2_132;
         pivot_in_2_133 <= pivot_out_2_132;
         start_in_2_133 <= start_out_2_132;
         swap_in_2_133 <= swap_out_2_132;
     end

     always @(posedge clk) begin
         data_in_2_133 <= data_out_1_133;
     end
  
     processor_AB AB_2_133 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_133),
       .start_in   (start_in_2_133),
       .swap_in   (swap_in_2_133),
       .op_in      (op_in_2_133),
       .pivot_in   (pivot_in_2_133),
       .start_out  (start_out_2_133),
       .swap_out   (swap_out_2_133),
       .data_out   (data_out_2_133),
       .op_out     (op_out_2_133),
       .pivot_out  (pivot_out_2_133),
       .r          (r_2_133)
     );

  // row 2, col 134

     reg start_in_2_134;
     wire start_out_2_134;

     reg swap_in_2_134;
     wire swap_out_2_134;

     reg [1:0] op_in_2_134;
     wire [1:0] op_out_2_134;

     wire r_2_134;

     reg data_in_2_134;
     wire data_out_2_134;

     reg pivot_in_2_134;
     wire pivot_out_2_134;

     always @(posedge clk) begin
         op_in_2_134 <= op_out_2_133;
         pivot_in_2_134 <= pivot_out_2_133;
         start_in_2_134 <= start_out_2_133;
         swap_in_2_134 <= swap_out_2_133;
     end

     always @(posedge clk) begin
         data_in_2_134 <= data_out_1_134;
     end
  
     processor_AB AB_2_134 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_134),
       .start_in   (start_in_2_134),
       .swap_in   (swap_in_2_134),
       .op_in      (op_in_2_134),
       .pivot_in   (pivot_in_2_134),
       .start_out  (start_out_2_134),
       .swap_out   (swap_out_2_134),
       .data_out   (data_out_2_134),
       .op_out     (op_out_2_134),
       .pivot_out  (pivot_out_2_134),
       .r          (r_2_134)
     );

  // row 2, col 135

     reg start_in_2_135;
     wire start_out_2_135;

     reg swap_in_2_135;
     wire swap_out_2_135;

     reg [1:0] op_in_2_135;
     wire [1:0] op_out_2_135;

     wire r_2_135;

     reg data_in_2_135;
     wire data_out_2_135;

     reg pivot_in_2_135;
     wire pivot_out_2_135;

     always @(posedge clk) begin
         op_in_2_135 <= op_out_2_134;
         pivot_in_2_135 <= pivot_out_2_134;
         start_in_2_135 <= start_out_2_134;
         swap_in_2_135 <= swap_out_2_134;
     end

     always @(posedge clk) begin
         data_in_2_135 <= data_out_1_135;
     end
  
     processor_AB AB_2_135 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_135),
       .start_in   (start_in_2_135),
       .swap_in   (swap_in_2_135),
       .op_in      (op_in_2_135),
       .pivot_in   (pivot_in_2_135),
       .start_out  (start_out_2_135),
       .swap_out   (swap_out_2_135),
       .data_out   (data_out_2_135),
       .op_out     (op_out_2_135),
       .pivot_out  (pivot_out_2_135),
       .r          (r_2_135)
     );

  // row 2, col 136

     reg start_in_2_136;
     wire start_out_2_136;

     reg swap_in_2_136;
     wire swap_out_2_136;

     reg [1:0] op_in_2_136;
     wire [1:0] op_out_2_136;

     wire r_2_136;

     reg data_in_2_136;
     wire data_out_2_136;

     reg pivot_in_2_136;
     wire pivot_out_2_136;

     always @(posedge clk) begin
         op_in_2_136 <= op_out_2_135;
         pivot_in_2_136 <= pivot_out_2_135;
         start_in_2_136 <= start_out_2_135;
         swap_in_2_136 <= swap_out_2_135;
     end

     always @(posedge clk) begin
         data_in_2_136 <= data_out_1_136;
     end
  
     processor_AB AB_2_136 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_136),
       .start_in   (start_in_2_136),
       .swap_in   (swap_in_2_136),
       .op_in      (op_in_2_136),
       .pivot_in   (pivot_in_2_136),
       .start_out  (start_out_2_136),
       .swap_out   (swap_out_2_136),
       .data_out   (data_out_2_136),
       .op_out     (op_out_2_136),
       .pivot_out  (pivot_out_2_136),
       .r          (r_2_136)
     );

  // row 2, col 137

     reg start_in_2_137;
     wire start_out_2_137;

     reg swap_in_2_137;
     wire swap_out_2_137;

     reg [1:0] op_in_2_137;
     wire [1:0] op_out_2_137;

     wire r_2_137;

     reg data_in_2_137;
     wire data_out_2_137;

     reg pivot_in_2_137;
     wire pivot_out_2_137;

     always @(posedge clk) begin
         op_in_2_137 <= op_out_2_136;
         pivot_in_2_137 <= pivot_out_2_136;
         start_in_2_137 <= start_out_2_136;
         swap_in_2_137 <= swap_out_2_136;
     end

     always @(posedge clk) begin
         data_in_2_137 <= data_out_1_137;
     end
  
     processor_AB AB_2_137 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_137),
       .start_in   (start_in_2_137),
       .swap_in   (swap_in_2_137),
       .op_in      (op_in_2_137),
       .pivot_in   (pivot_in_2_137),
       .start_out  (start_out_2_137),
       .swap_out   (swap_out_2_137),
       .data_out   (data_out_2_137),
       .op_out     (op_out_2_137),
       .pivot_out  (pivot_out_2_137),
       .r          (r_2_137)
     );

  // row 2, col 138

     reg start_in_2_138;
     wire start_out_2_138;

     reg swap_in_2_138;
     wire swap_out_2_138;

     reg [1:0] op_in_2_138;
     wire [1:0] op_out_2_138;

     wire r_2_138;

     reg data_in_2_138;
     wire data_out_2_138;

     reg pivot_in_2_138;
     wire pivot_out_2_138;

     always @(posedge clk) begin
         op_in_2_138 <= op_out_2_137;
         pivot_in_2_138 <= pivot_out_2_137;
         start_in_2_138 <= start_out_2_137;
         swap_in_2_138 <= swap_out_2_137;
     end

     always @(posedge clk) begin
         data_in_2_138 <= data_out_1_138;
     end
  
     processor_AB AB_2_138 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_138),
       .start_in   (start_in_2_138),
       .swap_in   (swap_in_2_138),
       .op_in      (op_in_2_138),
       .pivot_in   (pivot_in_2_138),
       .start_out  (start_out_2_138),
       .swap_out   (swap_out_2_138),
       .data_out   (data_out_2_138),
       .op_out     (op_out_2_138),
       .pivot_out  (pivot_out_2_138),
       .r          (r_2_138)
     );

  // row 2, col 139

     reg start_in_2_139;
     wire start_out_2_139;

     reg swap_in_2_139;
     wire swap_out_2_139;

     reg [1:0] op_in_2_139;
     wire [1:0] op_out_2_139;

     wire r_2_139;

     reg data_in_2_139;
     wire data_out_2_139;

     reg pivot_in_2_139;
     wire pivot_out_2_139;

     always @(posedge clk) begin
         op_in_2_139 <= op_out_2_138;
         pivot_in_2_139 <= pivot_out_2_138;
         start_in_2_139 <= start_out_2_138;
         swap_in_2_139 <= swap_out_2_138;
     end

     always @(posedge clk) begin
         data_in_2_139 <= data_out_1_139;
     end
  
     processor_AB AB_2_139 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_139),
       .start_in   (start_in_2_139),
       .swap_in   (swap_in_2_139),
       .op_in      (op_in_2_139),
       .pivot_in   (pivot_in_2_139),
       .start_out  (start_out_2_139),
       .swap_out   (swap_out_2_139),
       .data_out   (data_out_2_139),
       .op_out     (op_out_2_139),
       .pivot_out  (pivot_out_2_139),
       .r          (r_2_139)
     );

  // row 2, col 140

     reg start_in_2_140;
     wire start_out_2_140;

     reg swap_in_2_140;
     wire swap_out_2_140;

     reg [1:0] op_in_2_140;
     wire [1:0] op_out_2_140;

     wire r_2_140;

     reg data_in_2_140;
     wire data_out_2_140;

     reg pivot_in_2_140;
     wire pivot_out_2_140;

     always @(posedge clk) begin
         op_in_2_140 <= op_out_2_139;
         pivot_in_2_140 <= pivot_out_2_139;
         start_in_2_140 <= start_out_2_139;
         swap_in_2_140 <= swap_out_2_139;
     end

     always @(posedge clk) begin
         data_in_2_140 <= data_out_1_140;
     end
  
     processor_AB AB_2_140 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_140),
       .start_in   (start_in_2_140),
       .swap_in   (swap_in_2_140),
       .op_in      (op_in_2_140),
       .pivot_in   (pivot_in_2_140),
       .start_out  (start_out_2_140),
       .swap_out   (swap_out_2_140),
       .data_out   (data_out_2_140),
       .op_out     (op_out_2_140),
       .pivot_out  (pivot_out_2_140),
       .r          (r_2_140)
     );

  // row 2, col 141

     reg start_in_2_141;
     wire start_out_2_141;

     reg swap_in_2_141;
     wire swap_out_2_141;

     reg [1:0] op_in_2_141;
     wire [1:0] op_out_2_141;

     wire r_2_141;

     reg data_in_2_141;
     wire data_out_2_141;

     reg pivot_in_2_141;
     wire pivot_out_2_141;

     always @(posedge clk) begin
         op_in_2_141 <= op_out_2_140;
         pivot_in_2_141 <= pivot_out_2_140;
         start_in_2_141 <= start_out_2_140;
         swap_in_2_141 <= swap_out_2_140;
     end

     always @(posedge clk) begin
         data_in_2_141 <= data_out_1_141;
     end
  
     processor_AB AB_2_141 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_141),
       .start_in   (start_in_2_141),
       .swap_in   (swap_in_2_141),
       .op_in      (op_in_2_141),
       .pivot_in   (pivot_in_2_141),
       .start_out  (start_out_2_141),
       .swap_out   (swap_out_2_141),
       .data_out   (data_out_2_141),
       .op_out     (op_out_2_141),
       .pivot_out  (pivot_out_2_141),
       .r          (r_2_141)
     );

  // row 2, col 142

     reg start_in_2_142;
     wire start_out_2_142;

     reg swap_in_2_142;
     wire swap_out_2_142;

     reg [1:0] op_in_2_142;
     wire [1:0] op_out_2_142;

     wire r_2_142;

     reg data_in_2_142;
     wire data_out_2_142;

     reg pivot_in_2_142;
     wire pivot_out_2_142;

     always @(posedge clk) begin
         op_in_2_142 <= op_out_2_141;
         pivot_in_2_142 <= pivot_out_2_141;
         start_in_2_142 <= start_out_2_141;
         swap_in_2_142 <= swap_out_2_141;
     end

     always @(posedge clk) begin
         data_in_2_142 <= data_out_1_142;
     end
  
     processor_AB AB_2_142 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_142),
       .start_in   (start_in_2_142),
       .swap_in   (swap_in_2_142),
       .op_in      (op_in_2_142),
       .pivot_in   (pivot_in_2_142),
       .start_out  (start_out_2_142),
       .swap_out   (swap_out_2_142),
       .data_out   (data_out_2_142),
       .op_out     (op_out_2_142),
       .pivot_out  (pivot_out_2_142),
       .r          (r_2_142)
     );

  // row 2, col 143

     reg start_in_2_143;
     wire start_out_2_143;

     reg swap_in_2_143;
     wire swap_out_2_143;

     reg [1:0] op_in_2_143;
     wire [1:0] op_out_2_143;

     wire r_2_143;

     reg data_in_2_143;
     wire data_out_2_143;

     reg pivot_in_2_143;
     wire pivot_out_2_143;

     always @(posedge clk) begin
         op_in_2_143 <= op_out_2_142;
         pivot_in_2_143 <= pivot_out_2_142;
         start_in_2_143 <= start_out_2_142;
         swap_in_2_143 <= swap_out_2_142;
     end

     always @(posedge clk) begin
         data_in_2_143 <= data_out_1_143;
     end
  
     processor_AB AB_2_143 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_143),
       .start_in   (start_in_2_143),
       .swap_in   (swap_in_2_143),
       .op_in      (op_in_2_143),
       .pivot_in   (pivot_in_2_143),
       .start_out  (start_out_2_143),
       .swap_out   (swap_out_2_143),
       .data_out   (data_out_2_143),
       .op_out     (op_out_2_143),
       .pivot_out  (pivot_out_2_143),
       .r          (r_2_143)
     );

  // row 2, col 144

     reg start_in_2_144;
     wire start_out_2_144;

     reg swap_in_2_144;
     wire swap_out_2_144;

     reg [1:0] op_in_2_144;
     wire [1:0] op_out_2_144;

     wire r_2_144;

     reg data_in_2_144;
     wire data_out_2_144;

     reg pivot_in_2_144;
     wire pivot_out_2_144;

     always @(posedge clk) begin
         op_in_2_144 <= op_out_2_143;
         pivot_in_2_144 <= pivot_out_2_143;
         start_in_2_144 <= start_out_2_143;
         swap_in_2_144 <= swap_out_2_143;
     end

     always @(posedge clk) begin
         data_in_2_144 <= data_out_1_144;
     end
  
     processor_AB AB_2_144 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_144),
       .start_in   (start_in_2_144),
       .swap_in   (swap_in_2_144),
       .op_in      (op_in_2_144),
       .pivot_in   (pivot_in_2_144),
       .start_out  (start_out_2_144),
       .swap_out   (swap_out_2_144),
       .data_out   (data_out_2_144),
       .op_out     (op_out_2_144),
       .pivot_out  (pivot_out_2_144),
       .r          (r_2_144)
     );

  // row 2, col 145

     reg start_in_2_145;
     wire start_out_2_145;

     reg swap_in_2_145;
     wire swap_out_2_145;

     reg [1:0] op_in_2_145;
     wire [1:0] op_out_2_145;

     wire r_2_145;

     reg data_in_2_145;
     wire data_out_2_145;

     reg pivot_in_2_145;
     wire pivot_out_2_145;

     always @(posedge clk) begin
         op_in_2_145 <= op_out_2_144;
         pivot_in_2_145 <= pivot_out_2_144;
         start_in_2_145 <= start_out_2_144;
         swap_in_2_145 <= swap_out_2_144;
     end

     always @(posedge clk) begin
         data_in_2_145 <= data_out_1_145;
     end
  
     processor_AB AB_2_145 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_145),
       .start_in   (start_in_2_145),
       .swap_in   (swap_in_2_145),
       .op_in      (op_in_2_145),
       .pivot_in   (pivot_in_2_145),
       .start_out  (start_out_2_145),
       .swap_out   (swap_out_2_145),
       .data_out   (data_out_2_145),
       .op_out     (op_out_2_145),
       .pivot_out  (pivot_out_2_145),
       .r          (r_2_145)
     );

  // row 2, col 146

     reg start_in_2_146;
     wire start_out_2_146;

     reg swap_in_2_146;
     wire swap_out_2_146;

     reg [1:0] op_in_2_146;
     wire [1:0] op_out_2_146;

     wire r_2_146;

     reg data_in_2_146;
     wire data_out_2_146;

     reg pivot_in_2_146;
     wire pivot_out_2_146;

     always @(posedge clk) begin
         op_in_2_146 <= op_out_2_145;
         pivot_in_2_146 <= pivot_out_2_145;
         start_in_2_146 <= start_out_2_145;
         swap_in_2_146 <= swap_out_2_145;
     end

     always @(posedge clk) begin
         data_in_2_146 <= data_out_1_146;
     end
  
     processor_AB AB_2_146 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_146),
       .start_in   (start_in_2_146),
       .swap_in   (swap_in_2_146),
       .op_in      (op_in_2_146),
       .pivot_in   (pivot_in_2_146),
       .start_out  (start_out_2_146),
       .swap_out   (swap_out_2_146),
       .data_out   (data_out_2_146),
       .op_out     (op_out_2_146),
       .pivot_out  (pivot_out_2_146),
       .r          (r_2_146)
     );

  // row 2, col 147

     reg start_in_2_147;
     wire start_out_2_147;

     reg swap_in_2_147;
     wire swap_out_2_147;

     reg [1:0] op_in_2_147;
     wire [1:0] op_out_2_147;

     wire r_2_147;

     reg data_in_2_147;
     wire data_out_2_147;

     reg pivot_in_2_147;
     wire pivot_out_2_147;

     always @(posedge clk) begin
         op_in_2_147 <= op_out_2_146;
         pivot_in_2_147 <= pivot_out_2_146;
         start_in_2_147 <= start_out_2_146;
         swap_in_2_147 <= swap_out_2_146;
     end

     always @(posedge clk) begin
         data_in_2_147 <= data_out_1_147;
     end
  
     processor_AB AB_2_147 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_147),
       .start_in   (start_in_2_147),
       .swap_in   (swap_in_2_147),
       .op_in      (op_in_2_147),
       .pivot_in   (pivot_in_2_147),
       .start_out  (start_out_2_147),
       .swap_out   (swap_out_2_147),
       .data_out   (data_out_2_147),
       .op_out     (op_out_2_147),
       .pivot_out  (pivot_out_2_147),
       .r          (r_2_147)
     );

  // row 2, col 148

     reg start_in_2_148;
     wire start_out_2_148;

     reg swap_in_2_148;
     wire swap_out_2_148;

     reg [1:0] op_in_2_148;
     wire [1:0] op_out_2_148;

     wire r_2_148;

     reg data_in_2_148;
     wire data_out_2_148;

     reg pivot_in_2_148;
     wire pivot_out_2_148;

     always @(posedge clk) begin
         op_in_2_148 <= op_out_2_147;
         pivot_in_2_148 <= pivot_out_2_147;
         start_in_2_148 <= start_out_2_147;
         swap_in_2_148 <= swap_out_2_147;
     end

     always @(posedge clk) begin
         data_in_2_148 <= data_out_1_148;
     end
  
     processor_AB AB_2_148 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_148),
       .start_in   (start_in_2_148),
       .swap_in   (swap_in_2_148),
       .op_in      (op_in_2_148),
       .pivot_in   (pivot_in_2_148),
       .start_out  (start_out_2_148),
       .swap_out   (swap_out_2_148),
       .data_out   (data_out_2_148),
       .op_out     (op_out_2_148),
       .pivot_out  (pivot_out_2_148),
       .r          (r_2_148)
     );

  // row 2, col 149

     reg start_in_2_149;
     wire start_out_2_149;

     reg swap_in_2_149;
     wire swap_out_2_149;

     reg [1:0] op_in_2_149;
     wire [1:0] op_out_2_149;

     wire r_2_149;

     reg data_in_2_149;
     wire data_out_2_149;

     reg pivot_in_2_149;
     wire pivot_out_2_149;

     always @(posedge clk) begin
         op_in_2_149 <= op_out_2_148;
         pivot_in_2_149 <= pivot_out_2_148;
         start_in_2_149 <= start_out_2_148;
         swap_in_2_149 <= swap_out_2_148;
     end

     always @(posedge clk) begin
         data_in_2_149 <= data_out_1_149;
     end
  
     processor_AB AB_2_149 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_149),
       .start_in   (start_in_2_149),
       .swap_in   (swap_in_2_149),
       .op_in      (op_in_2_149),
       .pivot_in   (pivot_in_2_149),
       .start_out  (start_out_2_149),
       .swap_out   (swap_out_2_149),
       .data_out   (data_out_2_149),
       .op_out     (op_out_2_149),
       .pivot_out  (pivot_out_2_149),
       .r          (r_2_149)
     );

  // row 2, col 150

     reg start_in_2_150;
     wire start_out_2_150;

     reg swap_in_2_150;
     wire swap_out_2_150;

     reg [1:0] op_in_2_150;
     wire [1:0] op_out_2_150;

     wire r_2_150;

     reg data_in_2_150;
     wire data_out_2_150;

     reg pivot_in_2_150;
     wire pivot_out_2_150;

     always @(posedge clk) begin
         op_in_2_150 <= op_out_2_149;
         pivot_in_2_150 <= pivot_out_2_149;
         start_in_2_150 <= start_out_2_149;
         swap_in_2_150 <= swap_out_2_149;
     end

     always @(posedge clk) begin
         data_in_2_150 <= data_out_1_150;
     end
  
     processor_AB AB_2_150 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_150),
       .start_in   (start_in_2_150),
       .swap_in   (swap_in_2_150),
       .op_in      (op_in_2_150),
       .pivot_in   (pivot_in_2_150),
       .start_out  (start_out_2_150),
       .swap_out   (swap_out_2_150),
       .data_out   (data_out_2_150),
       .op_out     (op_out_2_150),
       .pivot_out  (pivot_out_2_150),
       .r          (r_2_150)
     );

  // row 2, col 151

     reg start_in_2_151;
     wire start_out_2_151;

     reg swap_in_2_151;
     wire swap_out_2_151;

     reg [1:0] op_in_2_151;
     wire [1:0] op_out_2_151;

     wire r_2_151;

     reg data_in_2_151;
     wire data_out_2_151;

     reg pivot_in_2_151;
     wire pivot_out_2_151;

     always @(posedge clk) begin
         op_in_2_151 <= op_out_2_150;
         pivot_in_2_151 <= pivot_out_2_150;
         start_in_2_151 <= start_out_2_150;
         swap_in_2_151 <= swap_out_2_150;
     end

     always @(posedge clk) begin
         data_in_2_151 <= data_out_1_151;
     end
  
     processor_AB AB_2_151 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_151),
       .start_in   (start_in_2_151),
       .swap_in   (swap_in_2_151),
       .op_in      (op_in_2_151),
       .pivot_in   (pivot_in_2_151),
       .start_out  (start_out_2_151),
       .swap_out   (swap_out_2_151),
       .data_out   (data_out_2_151),
       .op_out     (op_out_2_151),
       .pivot_out  (pivot_out_2_151),
       .r          (r_2_151)
     );

  // row 2, col 152

     reg start_in_2_152;
     wire start_out_2_152;

     reg swap_in_2_152;
     wire swap_out_2_152;

     reg [1:0] op_in_2_152;
     wire [1:0] op_out_2_152;

     wire r_2_152;

     reg data_in_2_152;
     wire data_out_2_152;

     reg pivot_in_2_152;
     wire pivot_out_2_152;

     always @(posedge clk) begin
         op_in_2_152 <= op_out_2_151;
         pivot_in_2_152 <= pivot_out_2_151;
         start_in_2_152 <= start_out_2_151;
         swap_in_2_152 <= swap_out_2_151;
     end

     always @(posedge clk) begin
         data_in_2_152 <= data_out_1_152;
     end
  
     processor_AB AB_2_152 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_152),
       .start_in   (start_in_2_152),
       .swap_in   (swap_in_2_152),
       .op_in      (op_in_2_152),
       .pivot_in   (pivot_in_2_152),
       .start_out  (start_out_2_152),
       .swap_out   (swap_out_2_152),
       .data_out   (data_out_2_152),
       .op_out     (op_out_2_152),
       .pivot_out  (pivot_out_2_152),
       .r          (r_2_152)
     );

  // row 2, col 153

     reg start_in_2_153;
     wire start_out_2_153;

     reg swap_in_2_153;
     wire swap_out_2_153;

     reg [1:0] op_in_2_153;
     wire [1:0] op_out_2_153;

     wire r_2_153;

     reg data_in_2_153;
     wire data_out_2_153;

     reg pivot_in_2_153;
     wire pivot_out_2_153;

     always @(posedge clk) begin
         op_in_2_153 <= op_out_2_152;
         pivot_in_2_153 <= pivot_out_2_152;
         start_in_2_153 <= start_out_2_152;
         swap_in_2_153 <= swap_out_2_152;
     end

     always @(posedge clk) begin
         data_in_2_153 <= data_out_1_153;
     end
  
     processor_AB AB_2_153 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_153),
       .start_in   (start_in_2_153),
       .swap_in   (swap_in_2_153),
       .op_in      (op_in_2_153),
       .pivot_in   (pivot_in_2_153),
       .start_out  (start_out_2_153),
       .swap_out   (swap_out_2_153),
       .data_out   (data_out_2_153),
       .op_out     (op_out_2_153),
       .pivot_out  (pivot_out_2_153),
       .r          (r_2_153)
     );

  // row 2, col 154

     reg start_in_2_154;
     wire start_out_2_154;

     reg swap_in_2_154;
     wire swap_out_2_154;

     reg [1:0] op_in_2_154;
     wire [1:0] op_out_2_154;

     wire r_2_154;

     reg data_in_2_154;
     wire data_out_2_154;

     reg pivot_in_2_154;
     wire pivot_out_2_154;

     always @(posedge clk) begin
         op_in_2_154 <= op_out_2_153;
         pivot_in_2_154 <= pivot_out_2_153;
         start_in_2_154 <= start_out_2_153;
         swap_in_2_154 <= swap_out_2_153;
     end

     always @(posedge clk) begin
         data_in_2_154 <= data_out_1_154;
     end
  
     processor_AB AB_2_154 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_154),
       .start_in   (start_in_2_154),
       .swap_in   (swap_in_2_154),
       .op_in      (op_in_2_154),
       .pivot_in   (pivot_in_2_154),
       .start_out  (start_out_2_154),
       .swap_out   (swap_out_2_154),
       .data_out   (data_out_2_154),
       .op_out     (op_out_2_154),
       .pivot_out  (pivot_out_2_154),
       .r          (r_2_154)
     );

  // row 2, col 155

     reg start_in_2_155;
     wire start_out_2_155;

     reg swap_in_2_155;
     wire swap_out_2_155;

     reg [1:0] op_in_2_155;
     wire [1:0] op_out_2_155;

     wire r_2_155;

     reg data_in_2_155;
     wire data_out_2_155;

     reg pivot_in_2_155;
     wire pivot_out_2_155;

     always @(posedge clk) begin
         op_in_2_155 <= op_out_2_154;
         pivot_in_2_155 <= pivot_out_2_154;
         start_in_2_155 <= start_out_2_154;
         swap_in_2_155 <= swap_out_2_154;
     end

     always @(posedge clk) begin
         data_in_2_155 <= data_out_1_155;
     end
  
     processor_AB AB_2_155 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_155),
       .start_in   (start_in_2_155),
       .swap_in   (swap_in_2_155),
       .op_in      (op_in_2_155),
       .pivot_in   (pivot_in_2_155),
       .start_out  (start_out_2_155),
       .swap_out   (swap_out_2_155),
       .data_out   (data_out_2_155),
       .op_out     (op_out_2_155),
       .pivot_out  (pivot_out_2_155),
       .r          (r_2_155)
     );

  // row 2, col 156

     reg start_in_2_156;
     wire start_out_2_156;

     reg swap_in_2_156;
     wire swap_out_2_156;

     reg [1:0] op_in_2_156;
     wire [1:0] op_out_2_156;

     wire r_2_156;

     reg data_in_2_156;
     wire data_out_2_156;

     reg pivot_in_2_156;
     wire pivot_out_2_156;

     always @(posedge clk) begin
         op_in_2_156 <= op_out_2_155;
         pivot_in_2_156 <= pivot_out_2_155;
         start_in_2_156 <= start_out_2_155;
         swap_in_2_156 <= swap_out_2_155;
     end

     always @(posedge clk) begin
         data_in_2_156 <= data_out_1_156;
     end
  
     processor_AB AB_2_156 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_156),
       .start_in   (start_in_2_156),
       .swap_in   (swap_in_2_156),
       .op_in      (op_in_2_156),
       .pivot_in   (pivot_in_2_156),
       .start_out  (start_out_2_156),
       .swap_out   (swap_out_2_156),
       .data_out   (data_out_2_156),
       .op_out     (op_out_2_156),
       .pivot_out  (pivot_out_2_156),
       .r          (r_2_156)
     );

  // row 2, col 157

     reg start_in_2_157;
     wire start_out_2_157;

     reg swap_in_2_157;
     wire swap_out_2_157;

     reg [1:0] op_in_2_157;
     wire [1:0] op_out_2_157;

     wire r_2_157;

     reg data_in_2_157;
     wire data_out_2_157;

     reg pivot_in_2_157;
     wire pivot_out_2_157;

     always @(posedge clk) begin
         op_in_2_157 <= op_out_2_156;
         pivot_in_2_157 <= pivot_out_2_156;
         start_in_2_157 <= start_out_2_156;
         swap_in_2_157 <= swap_out_2_156;
     end

     always @(posedge clk) begin
         data_in_2_157 <= data_out_1_157;
     end
  
     processor_AB AB_2_157 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_157),
       .start_in   (start_in_2_157),
       .swap_in   (swap_in_2_157),
       .op_in      (op_in_2_157),
       .pivot_in   (pivot_in_2_157),
       .start_out  (start_out_2_157),
       .swap_out   (swap_out_2_157),
       .data_out   (data_out_2_157),
       .op_out     (op_out_2_157),
       .pivot_out  (pivot_out_2_157),
       .r          (r_2_157)
     );

  // row 2, col 158

     reg start_in_2_158;
     wire start_out_2_158;

     reg swap_in_2_158;
     wire swap_out_2_158;

     reg [1:0] op_in_2_158;
     wire [1:0] op_out_2_158;

     wire r_2_158;

     reg data_in_2_158;
     wire data_out_2_158;

     reg pivot_in_2_158;
     wire pivot_out_2_158;

     always @(posedge clk) begin
         op_in_2_158 <= op_out_2_157;
         pivot_in_2_158 <= pivot_out_2_157;
         start_in_2_158 <= start_out_2_157;
         swap_in_2_158 <= swap_out_2_157;
     end

     always @(posedge clk) begin
         data_in_2_158 <= data_out_1_158;
     end
  
     processor_AB AB_2_158 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_158),
       .start_in   (start_in_2_158),
       .swap_in   (swap_in_2_158),
       .op_in      (op_in_2_158),
       .pivot_in   (pivot_in_2_158),
       .start_out  (start_out_2_158),
       .swap_out   (swap_out_2_158),
       .data_out   (data_out_2_158),
       .op_out     (op_out_2_158),
       .pivot_out  (pivot_out_2_158),
       .r          (r_2_158)
     );

  // row 2, col 159

     reg start_in_2_159;
     wire start_out_2_159;

     reg swap_in_2_159;
     wire swap_out_2_159;

     reg [1:0] op_in_2_159;
     wire [1:0] op_out_2_159;

     wire r_2_159;

     reg data_in_2_159;
     wire data_out_2_159;

     reg pivot_in_2_159;
     wire pivot_out_2_159;

     always @(posedge clk) begin
         op_in_2_159 <= op_out_2_158;
         pivot_in_2_159 <= pivot_out_2_158;
         start_in_2_159 <= start_out_2_158;
         swap_in_2_159 <= swap_out_2_158;
     end

     always @(posedge clk) begin
         data_in_2_159 <= data_out_1_159;
     end
  
     processor_AB AB_2_159 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_159),
       .start_in   (start_in_2_159),
       .swap_in   (swap_in_2_159),
       .op_in      (op_in_2_159),
       .pivot_in   (pivot_in_2_159),
       .start_out  (start_out_2_159),
       .swap_out   (swap_out_2_159),
       .data_out   (data_out_2_159),
       .op_out     (op_out_2_159),
       .pivot_out  (pivot_out_2_159),
       .r          (r_2_159)
     );

  // row 2, col 160

     reg start_in_2_160;
     wire start_out_2_160;

     reg swap_in_2_160;
     wire swap_out_2_160;

     reg [1:0] op_in_2_160;
     wire [1:0] op_out_2_160;

     wire r_2_160;

     reg data_in_2_160;
     wire data_out_2_160;

     reg pivot_in_2_160;
     wire pivot_out_2_160;

     always @(posedge clk) begin
         op_in_2_160 <= op_out_2_159;
         pivot_in_2_160 <= pivot_out_2_159;
         start_in_2_160 <= start_out_2_159;
         swap_in_2_160 <= swap_out_2_159;
     end

     always @(posedge clk) begin
         data_in_2_160 <= data_out_1_160;
     end
  
     processor_AB AB_2_160 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_160),
       .start_in   (start_in_2_160),
       .swap_in   (swap_in_2_160),
       .op_in      (op_in_2_160),
       .pivot_in   (pivot_in_2_160),
       .start_out  (start_out_2_160),
       .swap_out   (swap_out_2_160),
       .data_out   (data_out_2_160),
       .op_out     (op_out_2_160),
       .pivot_out  (pivot_out_2_160),
       .r          (r_2_160)
     );

  // row 2, col 161

     reg start_in_2_161;
     wire start_out_2_161;

     reg swap_in_2_161;
     wire swap_out_2_161;

     reg [1:0] op_in_2_161;
     wire [1:0] op_out_2_161;

     wire r_2_161;

     reg data_in_2_161;
     wire data_out_2_161;

     reg pivot_in_2_161;
     wire pivot_out_2_161;

     always @(posedge clk) begin
         op_in_2_161 <= op_out_2_160;
         pivot_in_2_161 <= pivot_out_2_160;
         start_in_2_161 <= start_out_2_160;
         swap_in_2_161 <= swap_out_2_160;
     end

     always @(posedge clk) begin
         data_in_2_161 <= data_out_1_161;
     end
  
     processor_AB AB_2_161 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_161),
       .start_in   (start_in_2_161),
       .swap_in   (swap_in_2_161),
       .op_in      (op_in_2_161),
       .pivot_in   (pivot_in_2_161),
       .start_out  (start_out_2_161),
       .swap_out   (swap_out_2_161),
       .data_out   (data_out_2_161),
       .op_out     (op_out_2_161),
       .pivot_out  (pivot_out_2_161),
       .r          (r_2_161)
     );

  // row 2, col 162

     reg start_in_2_162;
     wire start_out_2_162;

     reg swap_in_2_162;
     wire swap_out_2_162;

     reg [1:0] op_in_2_162;
     wire [1:0] op_out_2_162;

     wire r_2_162;

     reg data_in_2_162;
     wire data_out_2_162;

     reg pivot_in_2_162;
     wire pivot_out_2_162;

     always @(posedge clk) begin
         op_in_2_162 <= op_out_2_161;
         pivot_in_2_162 <= pivot_out_2_161;
         start_in_2_162 <= start_out_2_161;
         swap_in_2_162 <= swap_out_2_161;
     end

     always @(posedge clk) begin
         data_in_2_162 <= data_out_1_162;
     end
  
     processor_AB AB_2_162 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_162),
       .start_in   (start_in_2_162),
       .swap_in   (swap_in_2_162),
       .op_in      (op_in_2_162),
       .pivot_in   (pivot_in_2_162),
       .start_out  (start_out_2_162),
       .swap_out   (swap_out_2_162),
       .data_out   (data_out_2_162),
       .op_out     (op_out_2_162),
       .pivot_out  (pivot_out_2_162),
       .r          (r_2_162)
     );

  // row 2, col 163

     reg start_in_2_163;
     wire start_out_2_163;

     reg swap_in_2_163;
     wire swap_out_2_163;

     reg [1:0] op_in_2_163;
     wire [1:0] op_out_2_163;

     wire r_2_163;

     reg data_in_2_163;
     wire data_out_2_163;

     reg pivot_in_2_163;
     wire pivot_out_2_163;

     always @(posedge clk) begin
         op_in_2_163 <= op_out_2_162;
         pivot_in_2_163 <= pivot_out_2_162;
         start_in_2_163 <= start_out_2_162;
         swap_in_2_163 <= swap_out_2_162;
     end

     always @(posedge clk) begin
         data_in_2_163 <= data_out_1_163;
     end
  
     processor_AB AB_2_163 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_163),
       .start_in   (start_in_2_163),
       .swap_in   (swap_in_2_163),
       .op_in      (op_in_2_163),
       .pivot_in   (pivot_in_2_163),
       .start_out  (start_out_2_163),
       .swap_out   (swap_out_2_163),
       .data_out   (data_out_2_163),
       .op_out     (op_out_2_163),
       .pivot_out  (pivot_out_2_163),
       .r          (r_2_163)
     );

  // row 2, col 164

     reg start_in_2_164;
     wire start_out_2_164;

     reg swap_in_2_164;
     wire swap_out_2_164;

     reg [1:0] op_in_2_164;
     wire [1:0] op_out_2_164;

     wire r_2_164;

     reg data_in_2_164;
     wire data_out_2_164;

     reg pivot_in_2_164;
     wire pivot_out_2_164;

     always @(posedge clk) begin
         op_in_2_164 <= op_out_2_163;
         pivot_in_2_164 <= pivot_out_2_163;
         start_in_2_164 <= start_out_2_163;
         swap_in_2_164 <= swap_out_2_163;
     end

     always @(posedge clk) begin
         data_in_2_164 <= data_out_1_164;
     end
  
     processor_AB AB_2_164 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_164),
       .start_in   (start_in_2_164),
       .swap_in   (swap_in_2_164),
       .op_in      (op_in_2_164),
       .pivot_in   (pivot_in_2_164),
       .start_out  (start_out_2_164),
       .swap_out   (swap_out_2_164),
       .data_out   (data_out_2_164),
       .op_out     (op_out_2_164),
       .pivot_out  (pivot_out_2_164),
       .r          (r_2_164)
     );

  // row 2, col 165

     reg start_in_2_165;
     wire start_out_2_165;

     reg swap_in_2_165;
     wire swap_out_2_165;

     reg [1:0] op_in_2_165;
     wire [1:0] op_out_2_165;

     wire r_2_165;

     reg data_in_2_165;
     wire data_out_2_165;

     reg pivot_in_2_165;
     wire pivot_out_2_165;

     always @(posedge clk) begin
         op_in_2_165 <= op_out_2_164;
         pivot_in_2_165 <= pivot_out_2_164;
         start_in_2_165 <= start_out_2_164;
         swap_in_2_165 <= swap_out_2_164;
     end

     always @(posedge clk) begin
         data_in_2_165 <= data_out_1_165;
     end
  
     processor_AB AB_2_165 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_2_165),
       .start_in   (start_in_2_165),
       .swap_in   (swap_in_2_165),
       .op_in      (op_in_2_165),
       .pivot_in   (pivot_in_2_165),
       .start_out  (start_out_2_165),
       .swap_out   (swap_out_2_165),
       .data_out   (data_out_2_165),
       .op_out     (op_out_2_165),
       .pivot_out  (pivot_out_2_165),
       .r          (r_2_165)
     );

  /////////////////////////////////////
  // row 3
  // row 3, col 0

     wire start_in_3_0;
     wire start_out_3_0;

     wire swap_in_3_0;
     wire swap_out_3_0;

     wire [1:0] op_in_3_0;
     wire [1:0] op_out_3_0;

     wire r_3_0;

     reg data_in_3_0;
     wire data_out_3_0;

     wire pivot_in_3_0;
     wire pivout_out_3_0;

     assign op_in_3_0 = 2'b00;
     assign pivot_in_3_0 = 0;

     assign start_in_3_0 = start_row[3]; 
     assign swap_in_3_0 = mode ? swap : swap_row[3]; 

     always @(posedge clk) begin
         data_in_3_0 <= data_out_2_0;
     end

     processor_AB AB_3_0 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_0),
       .start_in   (start_in_3_0),
       .swap_in   (swap_in_3_0),
       .op_in      (op_in_3_0),
       .pivot_in   (pivot_in_3_0),
       .start_out  (start_out_3_0),
       .swap_out   (swap_out_3_0),
       .data_out   (data_out_3_0),
       .op_out     (op_out_3_0),
       .pivot_out  (pivot_out_3_0),
       .r          (r_3_0)
     );

  // row 3, col 1

     reg start_in_3_1;
     wire start_out_3_1;

     reg swap_in_3_1;
     wire swap_out_3_1;

     reg [1:0] op_in_3_1;
     wire [1:0] op_out_3_1;

     wire r_3_1;

     reg data_in_3_1;
     wire data_out_3_1;

     reg pivot_in_3_1;
     wire pivot_out_3_1;

     always @(posedge clk) begin
         op_in_3_1 <= op_out_3_0;
         pivot_in_3_1 <= pivot_out_3_0;
         start_in_3_1 <= start_out_3_0;
         swap_in_3_1 <= swap_out_3_0;
     end

     always @(posedge clk) begin
         data_in_3_1 <= data_out_2_1;
     end
  
     processor_AB AB_3_1 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_1),
       .start_in   (start_in_3_1),
       .swap_in   (swap_in_3_1),
       .op_in      (op_in_3_1),
       .pivot_in   (pivot_in_3_1),
       .start_out  (start_out_3_1),
       .swap_out   (swap_out_3_1),
       .data_out   (data_out_3_1),
       .op_out     (op_out_3_1),
       .pivot_out  (pivot_out_3_1),
       .r          (r_3_1)
     );

  // row 3, col 2

     reg start_in_3_2;
     wire start_out_3_2;

     reg swap_in_3_2;
     wire swap_out_3_2;

     reg [1:0] op_in_3_2;
     wire [1:0] op_out_3_2;

     wire r_3_2;

     reg data_in_3_2;
     wire data_out_3_2;

     reg pivot_in_3_2;
     wire pivot_out_3_2;

     always @(posedge clk) begin
         op_in_3_2 <= op_out_3_1;
         pivot_in_3_2 <= pivot_out_3_1;
         start_in_3_2 <= start_out_3_1;
         swap_in_3_2 <= swap_out_3_1;
     end

     always @(posedge clk) begin
         data_in_3_2 <= data_out_2_2;
     end
  
     processor_AB AB_3_2 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_2),
       .start_in   (start_in_3_2),
       .swap_in   (swap_in_3_2),
       .op_in      (op_in_3_2),
       .pivot_in   (pivot_in_3_2),
       .start_out  (start_out_3_2),
       .swap_out   (swap_out_3_2),
       .data_out   (data_out_3_2),
       .op_out     (op_out_3_2),
       .pivot_out  (pivot_out_3_2),
       .r          (r_3_2)
     );

  // row 3, col 3

     reg start_in_3_3;
     wire start_out_3_3;

     reg swap_in_3_3;
     wire swap_out_3_3;

     reg [1:0] op_in_3_3;
     wire [1:0] op_out_3_3;

     wire r_3_3;

     reg data_in_3_3;
     wire data_out_3_3;

     reg pivot_in_3_3;
     wire pivot_out_3_3;

     always @(posedge clk) begin
         op_in_3_3 <= op_out_3_2;
         pivot_in_3_3 <= pivot_out_3_2;
         start_in_3_3 <= start_out_3_2;
         swap_in_3_3 <= swap_out_3_2;
     end

     always @(posedge clk) begin
         data_in_3_3 <= data_out_2_3;
     end
  
     processor_AB AB_3_3 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_3),
       .start_in   (start_in_3_3),
       .swap_in   (swap_in_3_3),
       .op_in      (op_in_3_3),
       .pivot_in   (pivot_in_3_3),
       .start_out  (start_out_3_3),
       .swap_out   (swap_out_3_3),
       .data_out   (data_out_3_3),
       .op_out     (op_out_3_3),
       .pivot_out  (pivot_out_3_3),
       .r          (r_3_3)
     );

  // row 3, col 4

     reg start_in_3_4;
     wire start_out_3_4;

     reg swap_in_3_4;
     wire swap_out_3_4;

     reg [1:0] op_in_3_4;
     wire [1:0] op_out_3_4;

     wire r_3_4;

     reg data_in_3_4;
     wire data_out_3_4;

     reg pivot_in_3_4;
     wire pivot_out_3_4;

     always @(posedge clk) begin
         op_in_3_4 <= op_out_3_3;
         pivot_in_3_4 <= pivot_out_3_3;
         start_in_3_4 <= start_out_3_3;
         swap_in_3_4 <= swap_out_3_3;
     end

     always @(posedge clk) begin
         data_in_3_4 <= data_out_2_4;
     end
  
     processor_AB AB_3_4 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_4),
       .start_in   (start_in_3_4),
       .swap_in   (swap_in_3_4),
       .op_in      (op_in_3_4),
       .pivot_in   (pivot_in_3_4),
       .start_out  (start_out_3_4),
       .swap_out   (swap_out_3_4),
       .data_out   (data_out_3_4),
       .op_out     (op_out_3_4),
       .pivot_out  (pivot_out_3_4),
       .r          (r_3_4)
     );

  // row 3, col 5

     reg start_in_3_5;
     wire start_out_3_5;

     reg swap_in_3_5;
     wire swap_out_3_5;

     reg [1:0] op_in_3_5;
     wire [1:0] op_out_3_5;

     wire r_3_5;

     reg data_in_3_5;
     wire data_out_3_5;

     reg pivot_in_3_5;
     wire pivot_out_3_5;

     always @(posedge clk) begin
         op_in_3_5 <= op_out_3_4;
         pivot_in_3_5 <= pivot_out_3_4;
         start_in_3_5 <= start_out_3_4;
         swap_in_3_5 <= swap_out_3_4;
     end

     always @(posedge clk) begin
         data_in_3_5 <= data_out_2_5;
     end
  
     processor_AB AB_3_5 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_5),
       .start_in   (start_in_3_5),
       .swap_in   (swap_in_3_5),
       .op_in      (op_in_3_5),
       .pivot_in   (pivot_in_3_5),
       .start_out  (start_out_3_5),
       .swap_out   (swap_out_3_5),
       .data_out   (data_out_3_5),
       .op_out     (op_out_3_5),
       .pivot_out  (pivot_out_3_5),
       .r          (r_3_5)
     );

  // row 3, col 6

     reg start_in_3_6;
     wire start_out_3_6;

     reg swap_in_3_6;
     wire swap_out_3_6;

     reg [1:0] op_in_3_6;
     wire [1:0] op_out_3_6;

     wire r_3_6;

     reg data_in_3_6;
     wire data_out_3_6;

     reg pivot_in_3_6;
     wire pivot_out_3_6;

     always @(posedge clk) begin
         op_in_3_6 <= op_out_3_5;
         pivot_in_3_6 <= pivot_out_3_5;
         start_in_3_6 <= start_out_3_5;
         swap_in_3_6 <= swap_out_3_5;
     end

     always @(posedge clk) begin
         data_in_3_6 <= data_out_2_6;
     end
  
     processor_AB AB_3_6 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_6),
       .start_in   (start_in_3_6),
       .swap_in   (swap_in_3_6),
       .op_in      (op_in_3_6),
       .pivot_in   (pivot_in_3_6),
       .start_out  (start_out_3_6),
       .swap_out   (swap_out_3_6),
       .data_out   (data_out_3_6),
       .op_out     (op_out_3_6),
       .pivot_out  (pivot_out_3_6),
       .r          (r_3_6)
     );

  // row 3, col 7

     reg start_in_3_7;
     wire start_out_3_7;

     reg swap_in_3_7;
     wire swap_out_3_7;

     reg [1:0] op_in_3_7;
     wire [1:0] op_out_3_7;

     wire r_3_7;

     reg data_in_3_7;
     wire data_out_3_7;

     reg pivot_in_3_7;
     wire pivot_out_3_7;

     always @(posedge clk) begin
         op_in_3_7 <= op_out_3_6;
         pivot_in_3_7 <= pivot_out_3_6;
         start_in_3_7 <= start_out_3_6;
         swap_in_3_7 <= swap_out_3_6;
     end

     always @(posedge clk) begin
         data_in_3_7 <= data_out_2_7;
     end
  
     processor_AB AB_3_7 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_7),
       .start_in   (start_in_3_7),
       .swap_in   (swap_in_3_7),
       .op_in      (op_in_3_7),
       .pivot_in   (pivot_in_3_7),
       .start_out  (start_out_3_7),
       .swap_out   (swap_out_3_7),
       .data_out   (data_out_3_7),
       .op_out     (op_out_3_7),
       .pivot_out  (pivot_out_3_7),
       .r          (r_3_7)
     );

  // row 3, col 8

     reg start_in_3_8;
     wire start_out_3_8;

     reg swap_in_3_8;
     wire swap_out_3_8;

     reg [1:0] op_in_3_8;
     wire [1:0] op_out_3_8;

     wire r_3_8;

     reg data_in_3_8;
     wire data_out_3_8;

     reg pivot_in_3_8;
     wire pivot_out_3_8;

     always @(posedge clk) begin
         op_in_3_8 <= op_out_3_7;
         pivot_in_3_8 <= pivot_out_3_7;
         start_in_3_8 <= start_out_3_7;
         swap_in_3_8 <= swap_out_3_7;
     end

     always @(posedge clk) begin
         data_in_3_8 <= data_out_2_8;
     end
  
     processor_AB AB_3_8 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_8),
       .start_in   (start_in_3_8),
       .swap_in   (swap_in_3_8),
       .op_in      (op_in_3_8),
       .pivot_in   (pivot_in_3_8),
       .start_out  (start_out_3_8),
       .swap_out   (swap_out_3_8),
       .data_out   (data_out_3_8),
       .op_out     (op_out_3_8),
       .pivot_out  (pivot_out_3_8),
       .r          (r_3_8)
     );

  // row 3, col 9

     reg start_in_3_9;
     wire start_out_3_9;

     reg swap_in_3_9;
     wire swap_out_3_9;

     reg [1:0] op_in_3_9;
     wire [1:0] op_out_3_9;

     wire r_3_9;

     reg data_in_3_9;
     wire data_out_3_9;

     reg pivot_in_3_9;
     wire pivot_out_3_9;

     always @(posedge clk) begin
         op_in_3_9 <= op_out_3_8;
         pivot_in_3_9 <= pivot_out_3_8;
         start_in_3_9 <= start_out_3_8;
         swap_in_3_9 <= swap_out_3_8;
     end

     always @(posedge clk) begin
         data_in_3_9 <= data_out_2_9;
     end
  
     processor_AB AB_3_9 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_9),
       .start_in   (start_in_3_9),
       .swap_in   (swap_in_3_9),
       .op_in      (op_in_3_9),
       .pivot_in   (pivot_in_3_9),
       .start_out  (start_out_3_9),
       .swap_out   (swap_out_3_9),
       .data_out   (data_out_3_9),
       .op_out     (op_out_3_9),
       .pivot_out  (pivot_out_3_9),
       .r          (r_3_9)
     );

  // row 3, col 10

     reg start_in_3_10;
     wire start_out_3_10;

     reg swap_in_3_10;
     wire swap_out_3_10;

     reg [1:0] op_in_3_10;
     wire [1:0] op_out_3_10;

     wire r_3_10;

     reg data_in_3_10;
     wire data_out_3_10;

     reg pivot_in_3_10;
     wire pivot_out_3_10;

     always @(posedge clk) begin
         op_in_3_10 <= op_out_3_9;
         pivot_in_3_10 <= pivot_out_3_9;
         start_in_3_10 <= start_out_3_9;
         swap_in_3_10 <= swap_out_3_9;
     end

     always @(posedge clk) begin
         data_in_3_10 <= data_out_2_10;
     end
  
     processor_AB AB_3_10 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_10),
       .start_in   (start_in_3_10),
       .swap_in   (swap_in_3_10),
       .op_in      (op_in_3_10),
       .pivot_in   (pivot_in_3_10),
       .start_out  (start_out_3_10),
       .swap_out   (swap_out_3_10),
       .data_out   (data_out_3_10),
       .op_out     (op_out_3_10),
       .pivot_out  (pivot_out_3_10),
       .r          (r_3_10)
     );

  // row 3, col 11

     reg start_in_3_11;
     wire start_out_3_11;

     reg swap_in_3_11;
     wire swap_out_3_11;

     reg [1:0] op_in_3_11;
     wire [1:0] op_out_3_11;

     wire r_3_11;

     reg data_in_3_11;
     wire data_out_3_11;

     reg pivot_in_3_11;
     wire pivot_out_3_11;

     always @(posedge clk) begin
         op_in_3_11 <= op_out_3_10;
         pivot_in_3_11 <= pivot_out_3_10;
         start_in_3_11 <= start_out_3_10;
         swap_in_3_11 <= swap_out_3_10;
     end

     always @(posedge clk) begin
         data_in_3_11 <= data_out_2_11;
     end
  
     processor_AB AB_3_11 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_11),
       .start_in   (start_in_3_11),
       .swap_in   (swap_in_3_11),
       .op_in      (op_in_3_11),
       .pivot_in   (pivot_in_3_11),
       .start_out  (start_out_3_11),
       .swap_out   (swap_out_3_11),
       .data_out   (data_out_3_11),
       .op_out     (op_out_3_11),
       .pivot_out  (pivot_out_3_11),
       .r          (r_3_11)
     );

  // row 3, col 12

     reg start_in_3_12;
     wire start_out_3_12;

     reg swap_in_3_12;
     wire swap_out_3_12;

     reg [1:0] op_in_3_12;
     wire [1:0] op_out_3_12;

     wire r_3_12;

     reg data_in_3_12;
     wire data_out_3_12;

     reg pivot_in_3_12;
     wire pivot_out_3_12;

     always @(posedge clk) begin
         op_in_3_12 <= op_out_3_11;
         pivot_in_3_12 <= pivot_out_3_11;
         start_in_3_12 <= start_out_3_11;
         swap_in_3_12 <= swap_out_3_11;
     end

     always @(posedge clk) begin
         data_in_3_12 <= data_out_2_12;
     end
  
     processor_AB AB_3_12 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_12),
       .start_in   (start_in_3_12),
       .swap_in   (swap_in_3_12),
       .op_in      (op_in_3_12),
       .pivot_in   (pivot_in_3_12),
       .start_out  (start_out_3_12),
       .swap_out   (swap_out_3_12),
       .data_out   (data_out_3_12),
       .op_out     (op_out_3_12),
       .pivot_out  (pivot_out_3_12),
       .r          (r_3_12)
     );

  // row 3, col 13

     reg start_in_3_13;
     wire start_out_3_13;

     reg swap_in_3_13;
     wire swap_out_3_13;

     reg [1:0] op_in_3_13;
     wire [1:0] op_out_3_13;

     wire r_3_13;

     reg data_in_3_13;
     wire data_out_3_13;

     reg pivot_in_3_13;
     wire pivot_out_3_13;

     always @(posedge clk) begin
         op_in_3_13 <= op_out_3_12;
         pivot_in_3_13 <= pivot_out_3_12;
         start_in_3_13 <= start_out_3_12;
         swap_in_3_13 <= swap_out_3_12;
     end

     always @(posedge clk) begin
         data_in_3_13 <= data_out_2_13;
     end
  
     processor_AB AB_3_13 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_13),
       .start_in   (start_in_3_13),
       .swap_in   (swap_in_3_13),
       .op_in      (op_in_3_13),
       .pivot_in   (pivot_in_3_13),
       .start_out  (start_out_3_13),
       .swap_out   (swap_out_3_13),
       .data_out   (data_out_3_13),
       .op_out     (op_out_3_13),
       .pivot_out  (pivot_out_3_13),
       .r          (r_3_13)
     );

  // row 3, col 14

     reg start_in_3_14;
     wire start_out_3_14;

     reg swap_in_3_14;
     wire swap_out_3_14;

     reg [1:0] op_in_3_14;
     wire [1:0] op_out_3_14;

     wire r_3_14;

     reg data_in_3_14;
     wire data_out_3_14;

     reg pivot_in_3_14;
     wire pivot_out_3_14;

     always @(posedge clk) begin
         op_in_3_14 <= op_out_3_13;
         pivot_in_3_14 <= pivot_out_3_13;
         start_in_3_14 <= start_out_3_13;
         swap_in_3_14 <= swap_out_3_13;
     end

     always @(posedge clk) begin
         data_in_3_14 <= data_out_2_14;
     end
  
     processor_AB AB_3_14 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_14),
       .start_in   (start_in_3_14),
       .swap_in   (swap_in_3_14),
       .op_in      (op_in_3_14),
       .pivot_in   (pivot_in_3_14),
       .start_out  (start_out_3_14),
       .swap_out   (swap_out_3_14),
       .data_out   (data_out_3_14),
       .op_out     (op_out_3_14),
       .pivot_out  (pivot_out_3_14),
       .r          (r_3_14)
     );

  // row 3, col 15

     reg start_in_3_15;
     wire start_out_3_15;

     reg swap_in_3_15;
     wire swap_out_3_15;

     reg [1:0] op_in_3_15;
     wire [1:0] op_out_3_15;

     wire r_3_15;

     reg data_in_3_15;
     wire data_out_3_15;

     reg pivot_in_3_15;
     wire pivot_out_3_15;

     always @(posedge clk) begin
         op_in_3_15 <= op_out_3_14;
         pivot_in_3_15 <= pivot_out_3_14;
         start_in_3_15 <= start_out_3_14;
         swap_in_3_15 <= swap_out_3_14;
     end

     always @(posedge clk) begin
         data_in_3_15 <= data_out_2_15;
     end
  
     processor_AB AB_3_15 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_15),
       .start_in   (start_in_3_15),
       .swap_in   (swap_in_3_15),
       .op_in      (op_in_3_15),
       .pivot_in   (pivot_in_3_15),
       .start_out  (start_out_3_15),
       .swap_out   (swap_out_3_15),
       .data_out   (data_out_3_15),
       .op_out     (op_out_3_15),
       .pivot_out  (pivot_out_3_15),
       .r          (r_3_15)
     );

  // row 3, col 16

     reg start_in_3_16;
     wire start_out_3_16;

     reg swap_in_3_16;
     wire swap_out_3_16;

     reg [1:0] op_in_3_16;
     wire [1:0] op_out_3_16;

     wire r_3_16;

     reg data_in_3_16;
     wire data_out_3_16;

     reg pivot_in_3_16;
     wire pivot_out_3_16;

     always @(posedge clk) begin
         op_in_3_16 <= op_out_3_15;
         pivot_in_3_16 <= pivot_out_3_15;
         start_in_3_16 <= start_out_3_15;
         swap_in_3_16 <= swap_out_3_15;
     end

     always @(posedge clk) begin
         data_in_3_16 <= data_out_2_16;
     end
  
     processor_AB AB_3_16 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_16),
       .start_in   (start_in_3_16),
       .swap_in   (swap_in_3_16),
       .op_in      (op_in_3_16),
       .pivot_in   (pivot_in_3_16),
       .start_out  (start_out_3_16),
       .swap_out   (swap_out_3_16),
       .data_out   (data_out_3_16),
       .op_out     (op_out_3_16),
       .pivot_out  (pivot_out_3_16),
       .r          (r_3_16)
     );

  // row 3, col 17

     reg start_in_3_17;
     wire start_out_3_17;

     reg swap_in_3_17;
     wire swap_out_3_17;

     reg [1:0] op_in_3_17;
     wire [1:0] op_out_3_17;

     wire r_3_17;

     reg data_in_3_17;
     wire data_out_3_17;

     reg pivot_in_3_17;
     wire pivot_out_3_17;

     always @(posedge clk) begin
         op_in_3_17 <= op_out_3_16;
         pivot_in_3_17 <= pivot_out_3_16;
         start_in_3_17 <= start_out_3_16;
         swap_in_3_17 <= swap_out_3_16;
     end

     always @(posedge clk) begin
         data_in_3_17 <= data_out_2_17;
     end
  
     processor_AB AB_3_17 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_17),
       .start_in   (start_in_3_17),
       .swap_in   (swap_in_3_17),
       .op_in      (op_in_3_17),
       .pivot_in   (pivot_in_3_17),
       .start_out  (start_out_3_17),
       .swap_out   (swap_out_3_17),
       .data_out   (data_out_3_17),
       .op_out     (op_out_3_17),
       .pivot_out  (pivot_out_3_17),
       .r          (r_3_17)
     );

  // row 3, col 18

     reg start_in_3_18;
     wire start_out_3_18;

     reg swap_in_3_18;
     wire swap_out_3_18;

     reg [1:0] op_in_3_18;
     wire [1:0] op_out_3_18;

     wire r_3_18;

     reg data_in_3_18;
     wire data_out_3_18;

     reg pivot_in_3_18;
     wire pivot_out_3_18;

     always @(posedge clk) begin
         op_in_3_18 <= op_out_3_17;
         pivot_in_3_18 <= pivot_out_3_17;
         start_in_3_18 <= start_out_3_17;
         swap_in_3_18 <= swap_out_3_17;
     end

     always @(posedge clk) begin
         data_in_3_18 <= data_out_2_18;
     end
  
     processor_AB AB_3_18 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_18),
       .start_in   (start_in_3_18),
       .swap_in   (swap_in_3_18),
       .op_in      (op_in_3_18),
       .pivot_in   (pivot_in_3_18),
       .start_out  (start_out_3_18),
       .swap_out   (swap_out_3_18),
       .data_out   (data_out_3_18),
       .op_out     (op_out_3_18),
       .pivot_out  (pivot_out_3_18),
       .r          (r_3_18)
     );

  // row 3, col 19

     reg start_in_3_19;
     wire start_out_3_19;

     reg swap_in_3_19;
     wire swap_out_3_19;

     reg [1:0] op_in_3_19;
     wire [1:0] op_out_3_19;

     wire r_3_19;

     reg data_in_3_19;
     wire data_out_3_19;

     reg pivot_in_3_19;
     wire pivot_out_3_19;

     always @(posedge clk) begin
         op_in_3_19 <= op_out_3_18;
         pivot_in_3_19 <= pivot_out_3_18;
         start_in_3_19 <= start_out_3_18;
         swap_in_3_19 <= swap_out_3_18;
     end

     always @(posedge clk) begin
         data_in_3_19 <= data_out_2_19;
     end
  
     processor_AB AB_3_19 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_19),
       .start_in   (start_in_3_19),
       .swap_in   (swap_in_3_19),
       .op_in      (op_in_3_19),
       .pivot_in   (pivot_in_3_19),
       .start_out  (start_out_3_19),
       .swap_out   (swap_out_3_19),
       .data_out   (data_out_3_19),
       .op_out     (op_out_3_19),
       .pivot_out  (pivot_out_3_19),
       .r          (r_3_19)
     );

  // row 3, col 20

     reg start_in_3_20;
     wire start_out_3_20;

     reg swap_in_3_20;
     wire swap_out_3_20;

     reg [1:0] op_in_3_20;
     wire [1:0] op_out_3_20;

     wire r_3_20;

     reg data_in_3_20;
     wire data_out_3_20;

     reg pivot_in_3_20;
     wire pivot_out_3_20;

     always @(posedge clk) begin
         op_in_3_20 <= op_out_3_19;
         pivot_in_3_20 <= pivot_out_3_19;
         start_in_3_20 <= start_out_3_19;
         swap_in_3_20 <= swap_out_3_19;
     end

     always @(posedge clk) begin
         data_in_3_20 <= data_out_2_20;
     end
  
     processor_AB AB_3_20 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_20),
       .start_in   (start_in_3_20),
       .swap_in   (swap_in_3_20),
       .op_in      (op_in_3_20),
       .pivot_in   (pivot_in_3_20),
       .start_out  (start_out_3_20),
       .swap_out   (swap_out_3_20),
       .data_out   (data_out_3_20),
       .op_out     (op_out_3_20),
       .pivot_out  (pivot_out_3_20),
       .r          (r_3_20)
     );

  // row 3, col 21

     reg start_in_3_21;
     wire start_out_3_21;

     reg swap_in_3_21;
     wire swap_out_3_21;

     reg [1:0] op_in_3_21;
     wire [1:0] op_out_3_21;

     wire r_3_21;

     reg data_in_3_21;
     wire data_out_3_21;

     reg pivot_in_3_21;
     wire pivot_out_3_21;

     always @(posedge clk) begin
         op_in_3_21 <= op_out_3_20;
         pivot_in_3_21 <= pivot_out_3_20;
         start_in_3_21 <= start_out_3_20;
         swap_in_3_21 <= swap_out_3_20;
     end

     always @(posedge clk) begin
         data_in_3_21 <= data_out_2_21;
     end
  
     processor_AB AB_3_21 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_21),
       .start_in   (start_in_3_21),
       .swap_in   (swap_in_3_21),
       .op_in      (op_in_3_21),
       .pivot_in   (pivot_in_3_21),
       .start_out  (start_out_3_21),
       .swap_out   (swap_out_3_21),
       .data_out   (data_out_3_21),
       .op_out     (op_out_3_21),
       .pivot_out  (pivot_out_3_21),
       .r          (r_3_21)
     );

  // row 3, col 22

     reg start_in_3_22;
     wire start_out_3_22;

     reg swap_in_3_22;
     wire swap_out_3_22;

     reg [1:0] op_in_3_22;
     wire [1:0] op_out_3_22;

     wire r_3_22;

     reg data_in_3_22;
     wire data_out_3_22;

     reg pivot_in_3_22;
     wire pivot_out_3_22;

     always @(posedge clk) begin
         op_in_3_22 <= op_out_3_21;
         pivot_in_3_22 <= pivot_out_3_21;
         start_in_3_22 <= start_out_3_21;
         swap_in_3_22 <= swap_out_3_21;
     end

     always @(posedge clk) begin
         data_in_3_22 <= data_out_2_22;
     end
  
     processor_AB AB_3_22 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_22),
       .start_in   (start_in_3_22),
       .swap_in   (swap_in_3_22),
       .op_in      (op_in_3_22),
       .pivot_in   (pivot_in_3_22),
       .start_out  (start_out_3_22),
       .swap_out   (swap_out_3_22),
       .data_out   (data_out_3_22),
       .op_out     (op_out_3_22),
       .pivot_out  (pivot_out_3_22),
       .r          (r_3_22)
     );

  // row 3, col 23

     reg start_in_3_23;
     wire start_out_3_23;

     reg swap_in_3_23;
     wire swap_out_3_23;

     reg [1:0] op_in_3_23;
     wire [1:0] op_out_3_23;

     wire r_3_23;

     reg data_in_3_23;
     wire data_out_3_23;

     reg pivot_in_3_23;
     wire pivot_out_3_23;

     always @(posedge clk) begin
         op_in_3_23 <= op_out_3_22;
         pivot_in_3_23 <= pivot_out_3_22;
         start_in_3_23 <= start_out_3_22;
         swap_in_3_23 <= swap_out_3_22;
     end

     always @(posedge clk) begin
         data_in_3_23 <= data_out_2_23;
     end
  
     processor_AB AB_3_23 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_23),
       .start_in   (start_in_3_23),
       .swap_in   (swap_in_3_23),
       .op_in      (op_in_3_23),
       .pivot_in   (pivot_in_3_23),
       .start_out  (start_out_3_23),
       .swap_out   (swap_out_3_23),
       .data_out   (data_out_3_23),
       .op_out     (op_out_3_23),
       .pivot_out  (pivot_out_3_23),
       .r          (r_3_23)
     );

  // row 3, col 24

     reg start_in_3_24;
     wire start_out_3_24;

     reg swap_in_3_24;
     wire swap_out_3_24;

     reg [1:0] op_in_3_24;
     wire [1:0] op_out_3_24;

     wire r_3_24;

     reg data_in_3_24;
     wire data_out_3_24;

     reg pivot_in_3_24;
     wire pivot_out_3_24;

     always @(posedge clk) begin
         op_in_3_24 <= op_out_3_23;
         pivot_in_3_24 <= pivot_out_3_23;
         start_in_3_24 <= start_out_3_23;
         swap_in_3_24 <= swap_out_3_23;
     end

     always @(posedge clk) begin
         data_in_3_24 <= data_out_2_24;
     end
  
     processor_AB AB_3_24 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_24),
       .start_in   (start_in_3_24),
       .swap_in   (swap_in_3_24),
       .op_in      (op_in_3_24),
       .pivot_in   (pivot_in_3_24),
       .start_out  (start_out_3_24),
       .swap_out   (swap_out_3_24),
       .data_out   (data_out_3_24),
       .op_out     (op_out_3_24),
       .pivot_out  (pivot_out_3_24),
       .r          (r_3_24)
     );

  // row 3, col 25

     reg start_in_3_25;
     wire start_out_3_25;

     reg swap_in_3_25;
     wire swap_out_3_25;

     reg [1:0] op_in_3_25;
     wire [1:0] op_out_3_25;

     wire r_3_25;

     reg data_in_3_25;
     wire data_out_3_25;

     reg pivot_in_3_25;
     wire pivot_out_3_25;

     always @(posedge clk) begin
         op_in_3_25 <= op_out_3_24;
         pivot_in_3_25 <= pivot_out_3_24;
         start_in_3_25 <= start_out_3_24;
         swap_in_3_25 <= swap_out_3_24;
     end

     always @(posedge clk) begin
         data_in_3_25 <= data_out_2_25;
     end
  
     processor_AB AB_3_25 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_25),
       .start_in   (start_in_3_25),
       .swap_in   (swap_in_3_25),
       .op_in      (op_in_3_25),
       .pivot_in   (pivot_in_3_25),
       .start_out  (start_out_3_25),
       .swap_out   (swap_out_3_25),
       .data_out   (data_out_3_25),
       .op_out     (op_out_3_25),
       .pivot_out  (pivot_out_3_25),
       .r          (r_3_25)
     );

  // row 3, col 26

     reg start_in_3_26;
     wire start_out_3_26;

     reg swap_in_3_26;
     wire swap_out_3_26;

     reg [1:0] op_in_3_26;
     wire [1:0] op_out_3_26;

     wire r_3_26;

     reg data_in_3_26;
     wire data_out_3_26;

     reg pivot_in_3_26;
     wire pivot_out_3_26;

     always @(posedge clk) begin
         op_in_3_26 <= op_out_3_25;
         pivot_in_3_26 <= pivot_out_3_25;
         start_in_3_26 <= start_out_3_25;
         swap_in_3_26 <= swap_out_3_25;
     end

     always @(posedge clk) begin
         data_in_3_26 <= data_out_2_26;
     end
  
     processor_AB AB_3_26 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_26),
       .start_in   (start_in_3_26),
       .swap_in   (swap_in_3_26),
       .op_in      (op_in_3_26),
       .pivot_in   (pivot_in_3_26),
       .start_out  (start_out_3_26),
       .swap_out   (swap_out_3_26),
       .data_out   (data_out_3_26),
       .op_out     (op_out_3_26),
       .pivot_out  (pivot_out_3_26),
       .r          (r_3_26)
     );

  // row 3, col 27

     reg start_in_3_27;
     wire start_out_3_27;

     reg swap_in_3_27;
     wire swap_out_3_27;

     reg [1:0] op_in_3_27;
     wire [1:0] op_out_3_27;

     wire r_3_27;

     reg data_in_3_27;
     wire data_out_3_27;

     reg pivot_in_3_27;
     wire pivot_out_3_27;

     always @(posedge clk) begin
         op_in_3_27 <= op_out_3_26;
         pivot_in_3_27 <= pivot_out_3_26;
         start_in_3_27 <= start_out_3_26;
         swap_in_3_27 <= swap_out_3_26;
     end

     always @(posedge clk) begin
         data_in_3_27 <= data_out_2_27;
     end
  
     processor_AB AB_3_27 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_27),
       .start_in   (start_in_3_27),
       .swap_in   (swap_in_3_27),
       .op_in      (op_in_3_27),
       .pivot_in   (pivot_in_3_27),
       .start_out  (start_out_3_27),
       .swap_out   (swap_out_3_27),
       .data_out   (data_out_3_27),
       .op_out     (op_out_3_27),
       .pivot_out  (pivot_out_3_27),
       .r          (r_3_27)
     );

  // row 3, col 28

     reg start_in_3_28;
     wire start_out_3_28;

     reg swap_in_3_28;
     wire swap_out_3_28;

     reg [1:0] op_in_3_28;
     wire [1:0] op_out_3_28;

     wire r_3_28;

     reg data_in_3_28;
     wire data_out_3_28;

     reg pivot_in_3_28;
     wire pivot_out_3_28;

     always @(posedge clk) begin
         op_in_3_28 <= op_out_3_27;
         pivot_in_3_28 <= pivot_out_3_27;
         start_in_3_28 <= start_out_3_27;
         swap_in_3_28 <= swap_out_3_27;
     end

     always @(posedge clk) begin
         data_in_3_28 <= data_out_2_28;
     end
  
     processor_AB AB_3_28 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_28),
       .start_in   (start_in_3_28),
       .swap_in   (swap_in_3_28),
       .op_in      (op_in_3_28),
       .pivot_in   (pivot_in_3_28),
       .start_out  (start_out_3_28),
       .swap_out   (swap_out_3_28),
       .data_out   (data_out_3_28),
       .op_out     (op_out_3_28),
       .pivot_out  (pivot_out_3_28),
       .r          (r_3_28)
     );

  // row 3, col 29

     reg start_in_3_29;
     wire start_out_3_29;

     reg swap_in_3_29;
     wire swap_out_3_29;

     reg [1:0] op_in_3_29;
     wire [1:0] op_out_3_29;

     wire r_3_29;

     reg data_in_3_29;
     wire data_out_3_29;

     reg pivot_in_3_29;
     wire pivot_out_3_29;

     always @(posedge clk) begin
         op_in_3_29 <= op_out_3_28;
         pivot_in_3_29 <= pivot_out_3_28;
         start_in_3_29 <= start_out_3_28;
         swap_in_3_29 <= swap_out_3_28;
     end

     always @(posedge clk) begin
         data_in_3_29 <= data_out_2_29;
     end
  
     processor_AB AB_3_29 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_29),
       .start_in   (start_in_3_29),
       .swap_in   (swap_in_3_29),
       .op_in      (op_in_3_29),
       .pivot_in   (pivot_in_3_29),
       .start_out  (start_out_3_29),
       .swap_out   (swap_out_3_29),
       .data_out   (data_out_3_29),
       .op_out     (op_out_3_29),
       .pivot_out  (pivot_out_3_29),
       .r          (r_3_29)
     );

  // row 3, col 30

     reg start_in_3_30;
     wire start_out_3_30;

     reg swap_in_3_30;
     wire swap_out_3_30;

     reg [1:0] op_in_3_30;
     wire [1:0] op_out_3_30;

     wire r_3_30;

     reg data_in_3_30;
     wire data_out_3_30;

     reg pivot_in_3_30;
     wire pivot_out_3_30;

     always @(posedge clk) begin
         op_in_3_30 <= op_out_3_29;
         pivot_in_3_30 <= pivot_out_3_29;
         start_in_3_30 <= start_out_3_29;
         swap_in_3_30 <= swap_out_3_29;
     end

     always @(posedge clk) begin
         data_in_3_30 <= data_out_2_30;
     end
  
     processor_AB AB_3_30 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_30),
       .start_in   (start_in_3_30),
       .swap_in   (swap_in_3_30),
       .op_in      (op_in_3_30),
       .pivot_in   (pivot_in_3_30),
       .start_out  (start_out_3_30),
       .swap_out   (swap_out_3_30),
       .data_out   (data_out_3_30),
       .op_out     (op_out_3_30),
       .pivot_out  (pivot_out_3_30),
       .r          (r_3_30)
     );

  // row 3, col 31

     reg start_in_3_31;
     wire start_out_3_31;

     reg swap_in_3_31;
     wire swap_out_3_31;

     reg [1:0] op_in_3_31;
     wire [1:0] op_out_3_31;

     wire r_3_31;

     reg data_in_3_31;
     wire data_out_3_31;

     reg pivot_in_3_31;
     wire pivot_out_3_31;

     always @(posedge clk) begin
         op_in_3_31 <= op_out_3_30;
         pivot_in_3_31 <= pivot_out_3_30;
         start_in_3_31 <= start_out_3_30;
         swap_in_3_31 <= swap_out_3_30;
     end

     always @(posedge clk) begin
         data_in_3_31 <= data_out_2_31;
     end
  
     processor_AB AB_3_31 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_31),
       .start_in   (start_in_3_31),
       .swap_in   (swap_in_3_31),
       .op_in      (op_in_3_31),
       .pivot_in   (pivot_in_3_31),
       .start_out  (start_out_3_31),
       .swap_out   (swap_out_3_31),
       .data_out   (data_out_3_31),
       .op_out     (op_out_3_31),
       .pivot_out  (pivot_out_3_31),
       .r          (r_3_31)
     );

  // row 3, col 32

     reg start_in_3_32;
     wire start_out_3_32;

     reg swap_in_3_32;
     wire swap_out_3_32;

     reg [1:0] op_in_3_32;
     wire [1:0] op_out_3_32;

     wire r_3_32;

     reg data_in_3_32;
     wire data_out_3_32;

     reg pivot_in_3_32;
     wire pivot_out_3_32;

     always @(posedge clk) begin
         op_in_3_32 <= op_out_3_31;
         pivot_in_3_32 <= pivot_out_3_31;
         start_in_3_32 <= start_out_3_31;
         swap_in_3_32 <= swap_out_3_31;
     end

     always @(posedge clk) begin
         data_in_3_32 <= data_out_2_32;
     end
  
     processor_AB AB_3_32 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_32),
       .start_in   (start_in_3_32),
       .swap_in   (swap_in_3_32),
       .op_in      (op_in_3_32),
       .pivot_in   (pivot_in_3_32),
       .start_out  (start_out_3_32),
       .swap_out   (swap_out_3_32),
       .data_out   (data_out_3_32),
       .op_out     (op_out_3_32),
       .pivot_out  (pivot_out_3_32),
       .r          (r_3_32)
     );

  // row 3, col 33

     reg start_in_3_33;
     wire start_out_3_33;

     reg swap_in_3_33;
     wire swap_out_3_33;

     reg [1:0] op_in_3_33;
     wire [1:0] op_out_3_33;

     wire r_3_33;

     reg data_in_3_33;
     wire data_out_3_33;

     reg pivot_in_3_33;
     wire pivot_out_3_33;

     always @(posedge clk) begin
         op_in_3_33 <= op_out_3_32;
         pivot_in_3_33 <= pivot_out_3_32;
         start_in_3_33 <= start_out_3_32;
         swap_in_3_33 <= swap_out_3_32;
     end

     always @(posedge clk) begin
         data_in_3_33 <= data_out_2_33;
     end
  
     processor_AB AB_3_33 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_33),
       .start_in   (start_in_3_33),
       .swap_in   (swap_in_3_33),
       .op_in      (op_in_3_33),
       .pivot_in   (pivot_in_3_33),
       .start_out  (start_out_3_33),
       .swap_out   (swap_out_3_33),
       .data_out   (data_out_3_33),
       .op_out     (op_out_3_33),
       .pivot_out  (pivot_out_3_33),
       .r          (r_3_33)
     );

  // row 3, col 34

     reg start_in_3_34;
     wire start_out_3_34;

     reg swap_in_3_34;
     wire swap_out_3_34;

     reg [1:0] op_in_3_34;
     wire [1:0] op_out_3_34;

     wire r_3_34;

     reg data_in_3_34;
     wire data_out_3_34;

     reg pivot_in_3_34;
     wire pivot_out_3_34;

     always @(posedge clk) begin
         op_in_3_34 <= op_out_3_33;
         pivot_in_3_34 <= pivot_out_3_33;
         start_in_3_34 <= start_out_3_33;
         swap_in_3_34 <= swap_out_3_33;
     end

     always @(posedge clk) begin
         data_in_3_34 <= data_out_2_34;
     end
  
     processor_AB AB_3_34 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_34),
       .start_in   (start_in_3_34),
       .swap_in   (swap_in_3_34),
       .op_in      (op_in_3_34),
       .pivot_in   (pivot_in_3_34),
       .start_out  (start_out_3_34),
       .swap_out   (swap_out_3_34),
       .data_out   (data_out_3_34),
       .op_out     (op_out_3_34),
       .pivot_out  (pivot_out_3_34),
       .r          (r_3_34)
     );

  // row 3, col 35

     reg start_in_3_35;
     wire start_out_3_35;

     reg swap_in_3_35;
     wire swap_out_3_35;

     reg [1:0] op_in_3_35;
     wire [1:0] op_out_3_35;

     wire r_3_35;

     reg data_in_3_35;
     wire data_out_3_35;

     reg pivot_in_3_35;
     wire pivot_out_3_35;

     always @(posedge clk) begin
         op_in_3_35 <= op_out_3_34;
         pivot_in_3_35 <= pivot_out_3_34;
         start_in_3_35 <= start_out_3_34;
         swap_in_3_35 <= swap_out_3_34;
     end

     always @(posedge clk) begin
         data_in_3_35 <= data_out_2_35;
     end
  
     processor_AB AB_3_35 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_35),
       .start_in   (start_in_3_35),
       .swap_in   (swap_in_3_35),
       .op_in      (op_in_3_35),
       .pivot_in   (pivot_in_3_35),
       .start_out  (start_out_3_35),
       .swap_out   (swap_out_3_35),
       .data_out   (data_out_3_35),
       .op_out     (op_out_3_35),
       .pivot_out  (pivot_out_3_35),
       .r          (r_3_35)
     );

  // row 3, col 36

     reg start_in_3_36;
     wire start_out_3_36;

     reg swap_in_3_36;
     wire swap_out_3_36;

     reg [1:0] op_in_3_36;
     wire [1:0] op_out_3_36;

     wire r_3_36;

     reg data_in_3_36;
     wire data_out_3_36;

     reg pivot_in_3_36;
     wire pivot_out_3_36;

     always @(posedge clk) begin
         op_in_3_36 <= op_out_3_35;
         pivot_in_3_36 <= pivot_out_3_35;
         start_in_3_36 <= start_out_3_35;
         swap_in_3_36 <= swap_out_3_35;
     end

     always @(posedge clk) begin
         data_in_3_36 <= data_out_2_36;
     end
  
     processor_AB AB_3_36 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_36),
       .start_in   (start_in_3_36),
       .swap_in   (swap_in_3_36),
       .op_in      (op_in_3_36),
       .pivot_in   (pivot_in_3_36),
       .start_out  (start_out_3_36),
       .swap_out   (swap_out_3_36),
       .data_out   (data_out_3_36),
       .op_out     (op_out_3_36),
       .pivot_out  (pivot_out_3_36),
       .r          (r_3_36)
     );

  // row 3, col 37

     reg start_in_3_37;
     wire start_out_3_37;

     reg swap_in_3_37;
     wire swap_out_3_37;

     reg [1:0] op_in_3_37;
     wire [1:0] op_out_3_37;

     wire r_3_37;

     reg data_in_3_37;
     wire data_out_3_37;

     reg pivot_in_3_37;
     wire pivot_out_3_37;

     always @(posedge clk) begin
         op_in_3_37 <= op_out_3_36;
         pivot_in_3_37 <= pivot_out_3_36;
         start_in_3_37 <= start_out_3_36;
         swap_in_3_37 <= swap_out_3_36;
     end

     always @(posedge clk) begin
         data_in_3_37 <= data_out_2_37;
     end
  
     processor_AB AB_3_37 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_37),
       .start_in   (start_in_3_37),
       .swap_in   (swap_in_3_37),
       .op_in      (op_in_3_37),
       .pivot_in   (pivot_in_3_37),
       .start_out  (start_out_3_37),
       .swap_out   (swap_out_3_37),
       .data_out   (data_out_3_37),
       .op_out     (op_out_3_37),
       .pivot_out  (pivot_out_3_37),
       .r          (r_3_37)
     );

  // row 3, col 38

     reg start_in_3_38;
     wire start_out_3_38;

     reg swap_in_3_38;
     wire swap_out_3_38;

     reg [1:0] op_in_3_38;
     wire [1:0] op_out_3_38;

     wire r_3_38;

     reg data_in_3_38;
     wire data_out_3_38;

     reg pivot_in_3_38;
     wire pivot_out_3_38;

     always @(posedge clk) begin
         op_in_3_38 <= op_out_3_37;
         pivot_in_3_38 <= pivot_out_3_37;
         start_in_3_38 <= start_out_3_37;
         swap_in_3_38 <= swap_out_3_37;
     end

     always @(posedge clk) begin
         data_in_3_38 <= data_out_2_38;
     end
  
     processor_AB AB_3_38 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_38),
       .start_in   (start_in_3_38),
       .swap_in   (swap_in_3_38),
       .op_in      (op_in_3_38),
       .pivot_in   (pivot_in_3_38),
       .start_out  (start_out_3_38),
       .swap_out   (swap_out_3_38),
       .data_out   (data_out_3_38),
       .op_out     (op_out_3_38),
       .pivot_out  (pivot_out_3_38),
       .r          (r_3_38)
     );

  // row 3, col 39

     reg start_in_3_39;
     wire start_out_3_39;

     reg swap_in_3_39;
     wire swap_out_3_39;

     reg [1:0] op_in_3_39;
     wire [1:0] op_out_3_39;

     wire r_3_39;

     reg data_in_3_39;
     wire data_out_3_39;

     reg pivot_in_3_39;
     wire pivot_out_3_39;

     always @(posedge clk) begin
         op_in_3_39 <= op_out_3_38;
         pivot_in_3_39 <= pivot_out_3_38;
         start_in_3_39 <= start_out_3_38;
         swap_in_3_39 <= swap_out_3_38;
     end

     always @(posedge clk) begin
         data_in_3_39 <= data_out_2_39;
     end
  
     processor_AB AB_3_39 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_39),
       .start_in   (start_in_3_39),
       .swap_in   (swap_in_3_39),
       .op_in      (op_in_3_39),
       .pivot_in   (pivot_in_3_39),
       .start_out  (start_out_3_39),
       .swap_out   (swap_out_3_39),
       .data_out   (data_out_3_39),
       .op_out     (op_out_3_39),
       .pivot_out  (pivot_out_3_39),
       .r          (r_3_39)
     );

  // row 3, col 40

     reg start_in_3_40;
     wire start_out_3_40;

     reg swap_in_3_40;
     wire swap_out_3_40;

     reg [1:0] op_in_3_40;
     wire [1:0] op_out_3_40;

     wire r_3_40;

     reg data_in_3_40;
     wire data_out_3_40;

     reg pivot_in_3_40;
     wire pivot_out_3_40;

     always @(posedge clk) begin
         op_in_3_40 <= op_out_3_39;
         pivot_in_3_40 <= pivot_out_3_39;
         start_in_3_40 <= start_out_3_39;
         swap_in_3_40 <= swap_out_3_39;
     end

     always @(posedge clk) begin
         data_in_3_40 <= data_out_2_40;
     end
  
     processor_AB AB_3_40 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_40),
       .start_in   (start_in_3_40),
       .swap_in   (swap_in_3_40),
       .op_in      (op_in_3_40),
       .pivot_in   (pivot_in_3_40),
       .start_out  (start_out_3_40),
       .swap_out   (swap_out_3_40),
       .data_out   (data_out_3_40),
       .op_out     (op_out_3_40),
       .pivot_out  (pivot_out_3_40),
       .r          (r_3_40)
     );

  // row 3, col 41

     reg start_in_3_41;
     wire start_out_3_41;

     reg swap_in_3_41;
     wire swap_out_3_41;

     reg [1:0] op_in_3_41;
     wire [1:0] op_out_3_41;

     wire r_3_41;

     reg data_in_3_41;
     wire data_out_3_41;

     reg pivot_in_3_41;
     wire pivot_out_3_41;

     always @(posedge clk) begin
         op_in_3_41 <= op_out_3_40;
         pivot_in_3_41 <= pivot_out_3_40;
         start_in_3_41 <= start_out_3_40;
         swap_in_3_41 <= swap_out_3_40;
     end

     always @(posedge clk) begin
         data_in_3_41 <= data_out_2_41;
     end
  
     processor_AB AB_3_41 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_41),
       .start_in   (start_in_3_41),
       .swap_in   (swap_in_3_41),
       .op_in      (op_in_3_41),
       .pivot_in   (pivot_in_3_41),
       .start_out  (start_out_3_41),
       .swap_out   (swap_out_3_41),
       .data_out   (data_out_3_41),
       .op_out     (op_out_3_41),
       .pivot_out  (pivot_out_3_41),
       .r          (r_3_41)
     );

  // row 3, col 42

     reg start_in_3_42;
     wire start_out_3_42;

     reg swap_in_3_42;
     wire swap_out_3_42;

     reg [1:0] op_in_3_42;
     wire [1:0] op_out_3_42;

     wire r_3_42;

     reg data_in_3_42;
     wire data_out_3_42;

     reg pivot_in_3_42;
     wire pivot_out_3_42;

     always @(posedge clk) begin
         op_in_3_42 <= op_out_3_41;
         pivot_in_3_42 <= pivot_out_3_41;
         start_in_3_42 <= start_out_3_41;
         swap_in_3_42 <= swap_out_3_41;
     end

     always @(posedge clk) begin
         data_in_3_42 <= data_out_2_42;
     end
  
     processor_AB AB_3_42 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_42),
       .start_in   (start_in_3_42),
       .swap_in   (swap_in_3_42),
       .op_in      (op_in_3_42),
       .pivot_in   (pivot_in_3_42),
       .start_out  (start_out_3_42),
       .swap_out   (swap_out_3_42),
       .data_out   (data_out_3_42),
       .op_out     (op_out_3_42),
       .pivot_out  (pivot_out_3_42),
       .r          (r_3_42)
     );

  // row 3, col 43

     reg start_in_3_43;
     wire start_out_3_43;

     reg swap_in_3_43;
     wire swap_out_3_43;

     reg [1:0] op_in_3_43;
     wire [1:0] op_out_3_43;

     wire r_3_43;

     reg data_in_3_43;
     wire data_out_3_43;

     reg pivot_in_3_43;
     wire pivot_out_3_43;

     always @(posedge clk) begin
         op_in_3_43 <= op_out_3_42;
         pivot_in_3_43 <= pivot_out_3_42;
         start_in_3_43 <= start_out_3_42;
         swap_in_3_43 <= swap_out_3_42;
     end

     always @(posedge clk) begin
         data_in_3_43 <= data_out_2_43;
     end
  
     processor_AB AB_3_43 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_43),
       .start_in   (start_in_3_43),
       .swap_in   (swap_in_3_43),
       .op_in      (op_in_3_43),
       .pivot_in   (pivot_in_3_43),
       .start_out  (start_out_3_43),
       .swap_out   (swap_out_3_43),
       .data_out   (data_out_3_43),
       .op_out     (op_out_3_43),
       .pivot_out  (pivot_out_3_43),
       .r          (r_3_43)
     );

  // row 3, col 44

     reg start_in_3_44;
     wire start_out_3_44;

     reg swap_in_3_44;
     wire swap_out_3_44;

     reg [1:0] op_in_3_44;
     wire [1:0] op_out_3_44;

     wire r_3_44;

     reg data_in_3_44;
     wire data_out_3_44;

     reg pivot_in_3_44;
     wire pivot_out_3_44;

     always @(posedge clk) begin
         op_in_3_44 <= op_out_3_43;
         pivot_in_3_44 <= pivot_out_3_43;
         start_in_3_44 <= start_out_3_43;
         swap_in_3_44 <= swap_out_3_43;
     end

     always @(posedge clk) begin
         data_in_3_44 <= data_out_2_44;
     end
  
     processor_AB AB_3_44 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_44),
       .start_in   (start_in_3_44),
       .swap_in   (swap_in_3_44),
       .op_in      (op_in_3_44),
       .pivot_in   (pivot_in_3_44),
       .start_out  (start_out_3_44),
       .swap_out   (swap_out_3_44),
       .data_out   (data_out_3_44),
       .op_out     (op_out_3_44),
       .pivot_out  (pivot_out_3_44),
       .r          (r_3_44)
     );

  // row 3, col 45

     reg start_in_3_45;
     wire start_out_3_45;

     reg swap_in_3_45;
     wire swap_out_3_45;

     reg [1:0] op_in_3_45;
     wire [1:0] op_out_3_45;

     wire r_3_45;

     reg data_in_3_45;
     wire data_out_3_45;

     reg pivot_in_3_45;
     wire pivot_out_3_45;

     always @(posedge clk) begin
         op_in_3_45 <= op_out_3_44;
         pivot_in_3_45 <= pivot_out_3_44;
         start_in_3_45 <= start_out_3_44;
         swap_in_3_45 <= swap_out_3_44;
     end

     always @(posedge clk) begin
         data_in_3_45 <= data_out_2_45;
     end
  
     processor_AB AB_3_45 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_45),
       .start_in   (start_in_3_45),
       .swap_in   (swap_in_3_45),
       .op_in      (op_in_3_45),
       .pivot_in   (pivot_in_3_45),
       .start_out  (start_out_3_45),
       .swap_out   (swap_out_3_45),
       .data_out   (data_out_3_45),
       .op_out     (op_out_3_45),
       .pivot_out  (pivot_out_3_45),
       .r          (r_3_45)
     );

  // row 3, col 46

     reg start_in_3_46;
     wire start_out_3_46;

     reg swap_in_3_46;
     wire swap_out_3_46;

     reg [1:0] op_in_3_46;
     wire [1:0] op_out_3_46;

     wire r_3_46;

     reg data_in_3_46;
     wire data_out_3_46;

     reg pivot_in_3_46;
     wire pivot_out_3_46;

     always @(posedge clk) begin
         op_in_3_46 <= op_out_3_45;
         pivot_in_3_46 <= pivot_out_3_45;
         start_in_3_46 <= start_out_3_45;
         swap_in_3_46 <= swap_out_3_45;
     end

     always @(posedge clk) begin
         data_in_3_46 <= data_out_2_46;
     end
  
     processor_AB AB_3_46 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_46),
       .start_in   (start_in_3_46),
       .swap_in   (swap_in_3_46),
       .op_in      (op_in_3_46),
       .pivot_in   (pivot_in_3_46),
       .start_out  (start_out_3_46),
       .swap_out   (swap_out_3_46),
       .data_out   (data_out_3_46),
       .op_out     (op_out_3_46),
       .pivot_out  (pivot_out_3_46),
       .r          (r_3_46)
     );

  // row 3, col 47

     reg start_in_3_47;
     wire start_out_3_47;

     reg swap_in_3_47;
     wire swap_out_3_47;

     reg [1:0] op_in_3_47;
     wire [1:0] op_out_3_47;

     wire r_3_47;

     reg data_in_3_47;
     wire data_out_3_47;

     reg pivot_in_3_47;
     wire pivot_out_3_47;

     always @(posedge clk) begin
         op_in_3_47 <= op_out_3_46;
         pivot_in_3_47 <= pivot_out_3_46;
         start_in_3_47 <= start_out_3_46;
         swap_in_3_47 <= swap_out_3_46;
     end

     always @(posedge clk) begin
         data_in_3_47 <= data_out_2_47;
     end
  
     processor_AB AB_3_47 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_47),
       .start_in   (start_in_3_47),
       .swap_in   (swap_in_3_47),
       .op_in      (op_in_3_47),
       .pivot_in   (pivot_in_3_47),
       .start_out  (start_out_3_47),
       .swap_out   (swap_out_3_47),
       .data_out   (data_out_3_47),
       .op_out     (op_out_3_47),
       .pivot_out  (pivot_out_3_47),
       .r          (r_3_47)
     );

  // row 3, col 48

     reg start_in_3_48;
     wire start_out_3_48;

     reg swap_in_3_48;
     wire swap_out_3_48;

     reg [1:0] op_in_3_48;
     wire [1:0] op_out_3_48;

     wire r_3_48;

     reg data_in_3_48;
     wire data_out_3_48;

     reg pivot_in_3_48;
     wire pivot_out_3_48;

     always @(posedge clk) begin
         op_in_3_48 <= op_out_3_47;
         pivot_in_3_48 <= pivot_out_3_47;
         start_in_3_48 <= start_out_3_47;
         swap_in_3_48 <= swap_out_3_47;
     end

     always @(posedge clk) begin
         data_in_3_48 <= data_out_2_48;
     end
  
     processor_AB AB_3_48 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_48),
       .start_in   (start_in_3_48),
       .swap_in   (swap_in_3_48),
       .op_in      (op_in_3_48),
       .pivot_in   (pivot_in_3_48),
       .start_out  (start_out_3_48),
       .swap_out   (swap_out_3_48),
       .data_out   (data_out_3_48),
       .op_out     (op_out_3_48),
       .pivot_out  (pivot_out_3_48),
       .r          (r_3_48)
     );

  // row 3, col 49

     reg start_in_3_49;
     wire start_out_3_49;

     reg swap_in_3_49;
     wire swap_out_3_49;

     reg [1:0] op_in_3_49;
     wire [1:0] op_out_3_49;

     wire r_3_49;

     reg data_in_3_49;
     wire data_out_3_49;

     reg pivot_in_3_49;
     wire pivot_out_3_49;

     always @(posedge clk) begin
         op_in_3_49 <= op_out_3_48;
         pivot_in_3_49 <= pivot_out_3_48;
         start_in_3_49 <= start_out_3_48;
         swap_in_3_49 <= swap_out_3_48;
     end

     always @(posedge clk) begin
         data_in_3_49 <= data_out_2_49;
     end
  
     processor_AB AB_3_49 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_49),
       .start_in   (start_in_3_49),
       .swap_in   (swap_in_3_49),
       .op_in      (op_in_3_49),
       .pivot_in   (pivot_in_3_49),
       .start_out  (start_out_3_49),
       .swap_out   (swap_out_3_49),
       .data_out   (data_out_3_49),
       .op_out     (op_out_3_49),
       .pivot_out  (pivot_out_3_49),
       .r          (r_3_49)
     );

  // row 3, col 50

     reg start_in_3_50;
     wire start_out_3_50;

     reg swap_in_3_50;
     wire swap_out_3_50;

     reg [1:0] op_in_3_50;
     wire [1:0] op_out_3_50;

     wire r_3_50;

     reg data_in_3_50;
     wire data_out_3_50;

     reg pivot_in_3_50;
     wire pivot_out_3_50;

     always @(posedge clk) begin
         op_in_3_50 <= op_out_3_49;
         pivot_in_3_50 <= pivot_out_3_49;
         start_in_3_50 <= start_out_3_49;
         swap_in_3_50 <= swap_out_3_49;
     end

     always @(posedge clk) begin
         data_in_3_50 <= data_out_2_50;
     end
  
     processor_AB AB_3_50 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_50),
       .start_in   (start_in_3_50),
       .swap_in   (swap_in_3_50),
       .op_in      (op_in_3_50),
       .pivot_in   (pivot_in_3_50),
       .start_out  (start_out_3_50),
       .swap_out   (swap_out_3_50),
       .data_out   (data_out_3_50),
       .op_out     (op_out_3_50),
       .pivot_out  (pivot_out_3_50),
       .r          (r_3_50)
     );

  // row 3, col 51

     reg start_in_3_51;
     wire start_out_3_51;

     reg swap_in_3_51;
     wire swap_out_3_51;

     reg [1:0] op_in_3_51;
     wire [1:0] op_out_3_51;

     wire r_3_51;

     reg data_in_3_51;
     wire data_out_3_51;

     reg pivot_in_3_51;
     wire pivot_out_3_51;

     always @(posedge clk) begin
         op_in_3_51 <= op_out_3_50;
         pivot_in_3_51 <= pivot_out_3_50;
         start_in_3_51 <= start_out_3_50;
         swap_in_3_51 <= swap_out_3_50;
     end

     always @(posedge clk) begin
         data_in_3_51 <= data_out_2_51;
     end
  
     processor_AB AB_3_51 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_51),
       .start_in   (start_in_3_51),
       .swap_in   (swap_in_3_51),
       .op_in      (op_in_3_51),
       .pivot_in   (pivot_in_3_51),
       .start_out  (start_out_3_51),
       .swap_out   (swap_out_3_51),
       .data_out   (data_out_3_51),
       .op_out     (op_out_3_51),
       .pivot_out  (pivot_out_3_51),
       .r          (r_3_51)
     );

  // row 3, col 52

     reg start_in_3_52;
     wire start_out_3_52;

     reg swap_in_3_52;
     wire swap_out_3_52;

     reg [1:0] op_in_3_52;
     wire [1:0] op_out_3_52;

     wire r_3_52;

     reg data_in_3_52;
     wire data_out_3_52;

     reg pivot_in_3_52;
     wire pivot_out_3_52;

     always @(posedge clk) begin
         op_in_3_52 <= op_out_3_51;
         pivot_in_3_52 <= pivot_out_3_51;
         start_in_3_52 <= start_out_3_51;
         swap_in_3_52 <= swap_out_3_51;
     end

     always @(posedge clk) begin
         data_in_3_52 <= data_out_2_52;
     end
  
     processor_AB AB_3_52 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_52),
       .start_in   (start_in_3_52),
       .swap_in   (swap_in_3_52),
       .op_in      (op_in_3_52),
       .pivot_in   (pivot_in_3_52),
       .start_out  (start_out_3_52),
       .swap_out   (swap_out_3_52),
       .data_out   (data_out_3_52),
       .op_out     (op_out_3_52),
       .pivot_out  (pivot_out_3_52),
       .r          (r_3_52)
     );

  // row 3, col 53

     reg start_in_3_53;
     wire start_out_3_53;

     reg swap_in_3_53;
     wire swap_out_3_53;

     reg [1:0] op_in_3_53;
     wire [1:0] op_out_3_53;

     wire r_3_53;

     reg data_in_3_53;
     wire data_out_3_53;

     reg pivot_in_3_53;
     wire pivot_out_3_53;

     always @(posedge clk) begin
         op_in_3_53 <= op_out_3_52;
         pivot_in_3_53 <= pivot_out_3_52;
         start_in_3_53 <= start_out_3_52;
         swap_in_3_53 <= swap_out_3_52;
     end

     always @(posedge clk) begin
         data_in_3_53 <= data_out_2_53;
     end
  
     processor_AB AB_3_53 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_53),
       .start_in   (start_in_3_53),
       .swap_in   (swap_in_3_53),
       .op_in      (op_in_3_53),
       .pivot_in   (pivot_in_3_53),
       .start_out  (start_out_3_53),
       .swap_out   (swap_out_3_53),
       .data_out   (data_out_3_53),
       .op_out     (op_out_3_53),
       .pivot_out  (pivot_out_3_53),
       .r          (r_3_53)
     );

  // row 3, col 54

     reg start_in_3_54;
     wire start_out_3_54;

     reg swap_in_3_54;
     wire swap_out_3_54;

     reg [1:0] op_in_3_54;
     wire [1:0] op_out_3_54;

     wire r_3_54;

     reg data_in_3_54;
     wire data_out_3_54;

     reg pivot_in_3_54;
     wire pivot_out_3_54;

     always @(posedge clk) begin
         op_in_3_54 <= op_out_3_53;
         pivot_in_3_54 <= pivot_out_3_53;
         start_in_3_54 <= start_out_3_53;
         swap_in_3_54 <= swap_out_3_53;
     end

     always @(posedge clk) begin
         data_in_3_54 <= data_out_2_54;
     end
  
     processor_AB AB_3_54 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_54),
       .start_in   (start_in_3_54),
       .swap_in   (swap_in_3_54),
       .op_in      (op_in_3_54),
       .pivot_in   (pivot_in_3_54),
       .start_out  (start_out_3_54),
       .swap_out   (swap_out_3_54),
       .data_out   (data_out_3_54),
       .op_out     (op_out_3_54),
       .pivot_out  (pivot_out_3_54),
       .r          (r_3_54)
     );

  // row 3, col 55

     reg start_in_3_55;
     wire start_out_3_55;

     reg swap_in_3_55;
     wire swap_out_3_55;

     reg [1:0] op_in_3_55;
     wire [1:0] op_out_3_55;

     wire r_3_55;

     reg data_in_3_55;
     wire data_out_3_55;

     reg pivot_in_3_55;
     wire pivot_out_3_55;

     always @(posedge clk) begin
         op_in_3_55 <= op_out_3_54;
         pivot_in_3_55 <= pivot_out_3_54;
         start_in_3_55 <= start_out_3_54;
         swap_in_3_55 <= swap_out_3_54;
     end

     always @(posedge clk) begin
         data_in_3_55 <= data_out_2_55;
     end
  
     processor_AB AB_3_55 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_55),
       .start_in   (start_in_3_55),
       .swap_in   (swap_in_3_55),
       .op_in      (op_in_3_55),
       .pivot_in   (pivot_in_3_55),
       .start_out  (start_out_3_55),
       .swap_out   (swap_out_3_55),
       .data_out   (data_out_3_55),
       .op_out     (op_out_3_55),
       .pivot_out  (pivot_out_3_55),
       .r          (r_3_55)
     );

  // row 3, col 56

     reg start_in_3_56;
     wire start_out_3_56;

     reg swap_in_3_56;
     wire swap_out_3_56;

     reg [1:0] op_in_3_56;
     wire [1:0] op_out_3_56;

     wire r_3_56;

     reg data_in_3_56;
     wire data_out_3_56;

     reg pivot_in_3_56;
     wire pivot_out_3_56;

     always @(posedge clk) begin
         op_in_3_56 <= op_out_3_55;
         pivot_in_3_56 <= pivot_out_3_55;
         start_in_3_56 <= start_out_3_55;
         swap_in_3_56 <= swap_out_3_55;
     end

     always @(posedge clk) begin
         data_in_3_56 <= data_out_2_56;
     end
  
     processor_AB AB_3_56 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_56),
       .start_in   (start_in_3_56),
       .swap_in   (swap_in_3_56),
       .op_in      (op_in_3_56),
       .pivot_in   (pivot_in_3_56),
       .start_out  (start_out_3_56),
       .swap_out   (swap_out_3_56),
       .data_out   (data_out_3_56),
       .op_out     (op_out_3_56),
       .pivot_out  (pivot_out_3_56),
       .r          (r_3_56)
     );

  // row 3, col 57

     reg start_in_3_57;
     wire start_out_3_57;

     reg swap_in_3_57;
     wire swap_out_3_57;

     reg [1:0] op_in_3_57;
     wire [1:0] op_out_3_57;

     wire r_3_57;

     reg data_in_3_57;
     wire data_out_3_57;

     reg pivot_in_3_57;
     wire pivot_out_3_57;

     always @(posedge clk) begin
         op_in_3_57 <= op_out_3_56;
         pivot_in_3_57 <= pivot_out_3_56;
         start_in_3_57 <= start_out_3_56;
         swap_in_3_57 <= swap_out_3_56;
     end

     always @(posedge clk) begin
         data_in_3_57 <= data_out_2_57;
     end
  
     processor_AB AB_3_57 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_57),
       .start_in   (start_in_3_57),
       .swap_in   (swap_in_3_57),
       .op_in      (op_in_3_57),
       .pivot_in   (pivot_in_3_57),
       .start_out  (start_out_3_57),
       .swap_out   (swap_out_3_57),
       .data_out   (data_out_3_57),
       .op_out     (op_out_3_57),
       .pivot_out  (pivot_out_3_57),
       .r          (r_3_57)
     );

  // row 3, col 58

     reg start_in_3_58;
     wire start_out_3_58;

     reg swap_in_3_58;
     wire swap_out_3_58;

     reg [1:0] op_in_3_58;
     wire [1:0] op_out_3_58;

     wire r_3_58;

     reg data_in_3_58;
     wire data_out_3_58;

     reg pivot_in_3_58;
     wire pivot_out_3_58;

     always @(posedge clk) begin
         op_in_3_58 <= op_out_3_57;
         pivot_in_3_58 <= pivot_out_3_57;
         start_in_3_58 <= start_out_3_57;
         swap_in_3_58 <= swap_out_3_57;
     end

     always @(posedge clk) begin
         data_in_3_58 <= data_out_2_58;
     end
  
     processor_AB AB_3_58 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_58),
       .start_in   (start_in_3_58),
       .swap_in   (swap_in_3_58),
       .op_in      (op_in_3_58),
       .pivot_in   (pivot_in_3_58),
       .start_out  (start_out_3_58),
       .swap_out   (swap_out_3_58),
       .data_out   (data_out_3_58),
       .op_out     (op_out_3_58),
       .pivot_out  (pivot_out_3_58),
       .r          (r_3_58)
     );

  // row 3, col 59

     reg start_in_3_59;
     wire start_out_3_59;

     reg swap_in_3_59;
     wire swap_out_3_59;

     reg [1:0] op_in_3_59;
     wire [1:0] op_out_3_59;

     wire r_3_59;

     reg data_in_3_59;
     wire data_out_3_59;

     reg pivot_in_3_59;
     wire pivot_out_3_59;

     always @(posedge clk) begin
         op_in_3_59 <= op_out_3_58;
         pivot_in_3_59 <= pivot_out_3_58;
         start_in_3_59 <= start_out_3_58;
         swap_in_3_59 <= swap_out_3_58;
     end

     always @(posedge clk) begin
         data_in_3_59 <= data_out_2_59;
     end
  
     processor_AB AB_3_59 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_59),
       .start_in   (start_in_3_59),
       .swap_in   (swap_in_3_59),
       .op_in      (op_in_3_59),
       .pivot_in   (pivot_in_3_59),
       .start_out  (start_out_3_59),
       .swap_out   (swap_out_3_59),
       .data_out   (data_out_3_59),
       .op_out     (op_out_3_59),
       .pivot_out  (pivot_out_3_59),
       .r          (r_3_59)
     );

  // row 3, col 60

     reg start_in_3_60;
     wire start_out_3_60;

     reg swap_in_3_60;
     wire swap_out_3_60;

     reg [1:0] op_in_3_60;
     wire [1:0] op_out_3_60;

     wire r_3_60;

     reg data_in_3_60;
     wire data_out_3_60;

     reg pivot_in_3_60;
     wire pivot_out_3_60;

     always @(posedge clk) begin
         op_in_3_60 <= op_out_3_59;
         pivot_in_3_60 <= pivot_out_3_59;
         start_in_3_60 <= start_out_3_59;
         swap_in_3_60 <= swap_out_3_59;
     end

     always @(posedge clk) begin
         data_in_3_60 <= data_out_2_60;
     end
  
     processor_AB AB_3_60 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_60),
       .start_in   (start_in_3_60),
       .swap_in   (swap_in_3_60),
       .op_in      (op_in_3_60),
       .pivot_in   (pivot_in_3_60),
       .start_out  (start_out_3_60),
       .swap_out   (swap_out_3_60),
       .data_out   (data_out_3_60),
       .op_out     (op_out_3_60),
       .pivot_out  (pivot_out_3_60),
       .r          (r_3_60)
     );

  // row 3, col 61

     reg start_in_3_61;
     wire start_out_3_61;

     reg swap_in_3_61;
     wire swap_out_3_61;

     reg [1:0] op_in_3_61;
     wire [1:0] op_out_3_61;

     wire r_3_61;

     reg data_in_3_61;
     wire data_out_3_61;

     reg pivot_in_3_61;
     wire pivot_out_3_61;

     always @(posedge clk) begin
         op_in_3_61 <= op_out_3_60;
         pivot_in_3_61 <= pivot_out_3_60;
         start_in_3_61 <= start_out_3_60;
         swap_in_3_61 <= swap_out_3_60;
     end

     always @(posedge clk) begin
         data_in_3_61 <= data_out_2_61;
     end
  
     processor_AB AB_3_61 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_61),
       .start_in   (start_in_3_61),
       .swap_in   (swap_in_3_61),
       .op_in      (op_in_3_61),
       .pivot_in   (pivot_in_3_61),
       .start_out  (start_out_3_61),
       .swap_out   (swap_out_3_61),
       .data_out   (data_out_3_61),
       .op_out     (op_out_3_61),
       .pivot_out  (pivot_out_3_61),
       .r          (r_3_61)
     );

  // row 3, col 62

     reg start_in_3_62;
     wire start_out_3_62;

     reg swap_in_3_62;
     wire swap_out_3_62;

     reg [1:0] op_in_3_62;
     wire [1:0] op_out_3_62;

     wire r_3_62;

     reg data_in_3_62;
     wire data_out_3_62;

     reg pivot_in_3_62;
     wire pivot_out_3_62;

     always @(posedge clk) begin
         op_in_3_62 <= op_out_3_61;
         pivot_in_3_62 <= pivot_out_3_61;
         start_in_3_62 <= start_out_3_61;
         swap_in_3_62 <= swap_out_3_61;
     end

     always @(posedge clk) begin
         data_in_3_62 <= data_out_2_62;
     end
  
     processor_AB AB_3_62 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_62),
       .start_in   (start_in_3_62),
       .swap_in   (swap_in_3_62),
       .op_in      (op_in_3_62),
       .pivot_in   (pivot_in_3_62),
       .start_out  (start_out_3_62),
       .swap_out   (swap_out_3_62),
       .data_out   (data_out_3_62),
       .op_out     (op_out_3_62),
       .pivot_out  (pivot_out_3_62),
       .r          (r_3_62)
     );

  // row 3, col 63

     reg start_in_3_63;
     wire start_out_3_63;

     reg swap_in_3_63;
     wire swap_out_3_63;

     reg [1:0] op_in_3_63;
     wire [1:0] op_out_3_63;

     wire r_3_63;

     reg data_in_3_63;
     wire data_out_3_63;

     reg pivot_in_3_63;
     wire pivot_out_3_63;

     always @(posedge clk) begin
         op_in_3_63 <= op_out_3_62;
         pivot_in_3_63 <= pivot_out_3_62;
         start_in_3_63 <= start_out_3_62;
         swap_in_3_63 <= swap_out_3_62;
     end

     always @(posedge clk) begin
         data_in_3_63 <= data_out_2_63;
     end
  
     processor_AB AB_3_63 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_63),
       .start_in   (start_in_3_63),
       .swap_in   (swap_in_3_63),
       .op_in      (op_in_3_63),
       .pivot_in   (pivot_in_3_63),
       .start_out  (start_out_3_63),
       .swap_out   (swap_out_3_63),
       .data_out   (data_out_3_63),
       .op_out     (op_out_3_63),
       .pivot_out  (pivot_out_3_63),
       .r          (r_3_63)
     );

  // row 3, col 64

     reg start_in_3_64;
     wire start_out_3_64;

     reg swap_in_3_64;
     wire swap_out_3_64;

     reg [1:0] op_in_3_64;
     wire [1:0] op_out_3_64;

     wire r_3_64;

     reg data_in_3_64;
     wire data_out_3_64;

     reg pivot_in_3_64;
     wire pivot_out_3_64;

     always @(posedge clk) begin
         op_in_3_64 <= op_out_3_63;
         pivot_in_3_64 <= pivot_out_3_63;
         start_in_3_64 <= start_out_3_63;
         swap_in_3_64 <= swap_out_3_63;
     end

     always @(posedge clk) begin
         data_in_3_64 <= data_out_2_64;
     end
  
     processor_AB AB_3_64 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_64),
       .start_in   (start_in_3_64),
       .swap_in   (swap_in_3_64),
       .op_in      (op_in_3_64),
       .pivot_in   (pivot_in_3_64),
       .start_out  (start_out_3_64),
       .swap_out   (swap_out_3_64),
       .data_out   (data_out_3_64),
       .op_out     (op_out_3_64),
       .pivot_out  (pivot_out_3_64),
       .r          (r_3_64)
     );

  // row 3, col 65

     reg start_in_3_65;
     wire start_out_3_65;

     reg swap_in_3_65;
     wire swap_out_3_65;

     reg [1:0] op_in_3_65;
     wire [1:0] op_out_3_65;

     wire r_3_65;

     reg data_in_3_65;
     wire data_out_3_65;

     reg pivot_in_3_65;
     wire pivot_out_3_65;

     always @(posedge clk) begin
         op_in_3_65 <= op_out_3_64;
         pivot_in_3_65 <= pivot_out_3_64;
         start_in_3_65 <= start_out_3_64;
         swap_in_3_65 <= swap_out_3_64;
     end

     always @(posedge clk) begin
         data_in_3_65 <= data_out_2_65;
     end
  
     processor_AB AB_3_65 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_65),
       .start_in   (start_in_3_65),
       .swap_in   (swap_in_3_65),
       .op_in      (op_in_3_65),
       .pivot_in   (pivot_in_3_65),
       .start_out  (start_out_3_65),
       .swap_out   (swap_out_3_65),
       .data_out   (data_out_3_65),
       .op_out     (op_out_3_65),
       .pivot_out  (pivot_out_3_65),
       .r          (r_3_65)
     );

  // row 3, col 66

     reg start_in_3_66;
     wire start_out_3_66;

     reg swap_in_3_66;
     wire swap_out_3_66;

     reg [1:0] op_in_3_66;
     wire [1:0] op_out_3_66;

     wire r_3_66;

     reg data_in_3_66;
     wire data_out_3_66;

     reg pivot_in_3_66;
     wire pivot_out_3_66;

     always @(posedge clk) begin
         op_in_3_66 <= op_out_3_65;
         pivot_in_3_66 <= pivot_out_3_65;
         start_in_3_66 <= start_out_3_65;
         swap_in_3_66 <= swap_out_3_65;
     end

     always @(posedge clk) begin
         data_in_3_66 <= data_out_2_66;
     end
  
     processor_AB AB_3_66 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_66),
       .start_in   (start_in_3_66),
       .swap_in   (swap_in_3_66),
       .op_in      (op_in_3_66),
       .pivot_in   (pivot_in_3_66),
       .start_out  (start_out_3_66),
       .swap_out   (swap_out_3_66),
       .data_out   (data_out_3_66),
       .op_out     (op_out_3_66),
       .pivot_out  (pivot_out_3_66),
       .r          (r_3_66)
     );

  // row 3, col 67

     reg start_in_3_67;
     wire start_out_3_67;

     reg swap_in_3_67;
     wire swap_out_3_67;

     reg [1:0] op_in_3_67;
     wire [1:0] op_out_3_67;

     wire r_3_67;

     reg data_in_3_67;
     wire data_out_3_67;

     reg pivot_in_3_67;
     wire pivot_out_3_67;

     always @(posedge clk) begin
         op_in_3_67 <= op_out_3_66;
         pivot_in_3_67 <= pivot_out_3_66;
         start_in_3_67 <= start_out_3_66;
         swap_in_3_67 <= swap_out_3_66;
     end

     always @(posedge clk) begin
         data_in_3_67 <= data_out_2_67;
     end
  
     processor_AB AB_3_67 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_67),
       .start_in   (start_in_3_67),
       .swap_in   (swap_in_3_67),
       .op_in      (op_in_3_67),
       .pivot_in   (pivot_in_3_67),
       .start_out  (start_out_3_67),
       .swap_out   (swap_out_3_67),
       .data_out   (data_out_3_67),
       .op_out     (op_out_3_67),
       .pivot_out  (pivot_out_3_67),
       .r          (r_3_67)
     );

  // row 3, col 68

     reg start_in_3_68;
     wire start_out_3_68;

     reg swap_in_3_68;
     wire swap_out_3_68;

     reg [1:0] op_in_3_68;
     wire [1:0] op_out_3_68;

     wire r_3_68;

     reg data_in_3_68;
     wire data_out_3_68;

     reg pivot_in_3_68;
     wire pivot_out_3_68;

     always @(posedge clk) begin
         op_in_3_68 <= op_out_3_67;
         pivot_in_3_68 <= pivot_out_3_67;
         start_in_3_68 <= start_out_3_67;
         swap_in_3_68 <= swap_out_3_67;
     end

     always @(posedge clk) begin
         data_in_3_68 <= data_out_2_68;
     end
  
     processor_AB AB_3_68 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_68),
       .start_in   (start_in_3_68),
       .swap_in   (swap_in_3_68),
       .op_in      (op_in_3_68),
       .pivot_in   (pivot_in_3_68),
       .start_out  (start_out_3_68),
       .swap_out   (swap_out_3_68),
       .data_out   (data_out_3_68),
       .op_out     (op_out_3_68),
       .pivot_out  (pivot_out_3_68),
       .r          (r_3_68)
     );

  // row 3, col 69

     reg start_in_3_69;
     wire start_out_3_69;

     reg swap_in_3_69;
     wire swap_out_3_69;

     reg [1:0] op_in_3_69;
     wire [1:0] op_out_3_69;

     wire r_3_69;

     reg data_in_3_69;
     wire data_out_3_69;

     reg pivot_in_3_69;
     wire pivot_out_3_69;

     always @(posedge clk) begin
         op_in_3_69 <= op_out_3_68;
         pivot_in_3_69 <= pivot_out_3_68;
         start_in_3_69 <= start_out_3_68;
         swap_in_3_69 <= swap_out_3_68;
     end

     always @(posedge clk) begin
         data_in_3_69 <= data_out_2_69;
     end
  
     processor_AB AB_3_69 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_69),
       .start_in   (start_in_3_69),
       .swap_in   (swap_in_3_69),
       .op_in      (op_in_3_69),
       .pivot_in   (pivot_in_3_69),
       .start_out  (start_out_3_69),
       .swap_out   (swap_out_3_69),
       .data_out   (data_out_3_69),
       .op_out     (op_out_3_69),
       .pivot_out  (pivot_out_3_69),
       .r          (r_3_69)
     );

  // row 3, col 70

     reg start_in_3_70;
     wire start_out_3_70;

     reg swap_in_3_70;
     wire swap_out_3_70;

     reg [1:0] op_in_3_70;
     wire [1:0] op_out_3_70;

     wire r_3_70;

     reg data_in_3_70;
     wire data_out_3_70;

     reg pivot_in_3_70;
     wire pivot_out_3_70;

     always @(posedge clk) begin
         op_in_3_70 <= op_out_3_69;
         pivot_in_3_70 <= pivot_out_3_69;
         start_in_3_70 <= start_out_3_69;
         swap_in_3_70 <= swap_out_3_69;
     end

     always @(posedge clk) begin
         data_in_3_70 <= data_out_2_70;
     end
  
     processor_AB AB_3_70 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_70),
       .start_in   (start_in_3_70),
       .swap_in   (swap_in_3_70),
       .op_in      (op_in_3_70),
       .pivot_in   (pivot_in_3_70),
       .start_out  (start_out_3_70),
       .swap_out   (swap_out_3_70),
       .data_out   (data_out_3_70),
       .op_out     (op_out_3_70),
       .pivot_out  (pivot_out_3_70),
       .r          (r_3_70)
     );

  // row 3, col 71

     reg start_in_3_71;
     wire start_out_3_71;

     reg swap_in_3_71;
     wire swap_out_3_71;

     reg [1:0] op_in_3_71;
     wire [1:0] op_out_3_71;

     wire r_3_71;

     reg data_in_3_71;
     wire data_out_3_71;

     reg pivot_in_3_71;
     wire pivot_out_3_71;

     always @(posedge clk) begin
         op_in_3_71 <= op_out_3_70;
         pivot_in_3_71 <= pivot_out_3_70;
         start_in_3_71 <= start_out_3_70;
         swap_in_3_71 <= swap_out_3_70;
     end

     always @(posedge clk) begin
         data_in_3_71 <= data_out_2_71;
     end
  
     processor_AB AB_3_71 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_71),
       .start_in   (start_in_3_71),
       .swap_in   (swap_in_3_71),
       .op_in      (op_in_3_71),
       .pivot_in   (pivot_in_3_71),
       .start_out  (start_out_3_71),
       .swap_out   (swap_out_3_71),
       .data_out   (data_out_3_71),
       .op_out     (op_out_3_71),
       .pivot_out  (pivot_out_3_71),
       .r          (r_3_71)
     );

  // row 3, col 72

     reg start_in_3_72;
     wire start_out_3_72;

     reg swap_in_3_72;
     wire swap_out_3_72;

     reg [1:0] op_in_3_72;
     wire [1:0] op_out_3_72;

     wire r_3_72;

     reg data_in_3_72;
     wire data_out_3_72;

     reg pivot_in_3_72;
     wire pivot_out_3_72;

     always @(posedge clk) begin
         op_in_3_72 <= op_out_3_71;
         pivot_in_3_72 <= pivot_out_3_71;
         start_in_3_72 <= start_out_3_71;
         swap_in_3_72 <= swap_out_3_71;
     end

     always @(posedge clk) begin
         data_in_3_72 <= data_out_2_72;
     end
  
     processor_AB AB_3_72 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_72),
       .start_in   (start_in_3_72),
       .swap_in   (swap_in_3_72),
       .op_in      (op_in_3_72),
       .pivot_in   (pivot_in_3_72),
       .start_out  (start_out_3_72),
       .swap_out   (swap_out_3_72),
       .data_out   (data_out_3_72),
       .op_out     (op_out_3_72),
       .pivot_out  (pivot_out_3_72),
       .r          (r_3_72)
     );

  // row 3, col 73

     reg start_in_3_73;
     wire start_out_3_73;

     reg swap_in_3_73;
     wire swap_out_3_73;

     reg [1:0] op_in_3_73;
     wire [1:0] op_out_3_73;

     wire r_3_73;

     reg data_in_3_73;
     wire data_out_3_73;

     reg pivot_in_3_73;
     wire pivot_out_3_73;

     always @(posedge clk) begin
         op_in_3_73 <= op_out_3_72;
         pivot_in_3_73 <= pivot_out_3_72;
         start_in_3_73 <= start_out_3_72;
         swap_in_3_73 <= swap_out_3_72;
     end

     always @(posedge clk) begin
         data_in_3_73 <= data_out_2_73;
     end
  
     processor_AB AB_3_73 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_73),
       .start_in   (start_in_3_73),
       .swap_in   (swap_in_3_73),
       .op_in      (op_in_3_73),
       .pivot_in   (pivot_in_3_73),
       .start_out  (start_out_3_73),
       .swap_out   (swap_out_3_73),
       .data_out   (data_out_3_73),
       .op_out     (op_out_3_73),
       .pivot_out  (pivot_out_3_73),
       .r          (r_3_73)
     );

  // row 3, col 74

     reg start_in_3_74;
     wire start_out_3_74;

     reg swap_in_3_74;
     wire swap_out_3_74;

     reg [1:0] op_in_3_74;
     wire [1:0] op_out_3_74;

     wire r_3_74;

     reg data_in_3_74;
     wire data_out_3_74;

     reg pivot_in_3_74;
     wire pivot_out_3_74;

     always @(posedge clk) begin
         op_in_3_74 <= op_out_3_73;
         pivot_in_3_74 <= pivot_out_3_73;
         start_in_3_74 <= start_out_3_73;
         swap_in_3_74 <= swap_out_3_73;
     end

     always @(posedge clk) begin
         data_in_3_74 <= data_out_2_74;
     end
  
     processor_AB AB_3_74 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_74),
       .start_in   (start_in_3_74),
       .swap_in   (swap_in_3_74),
       .op_in      (op_in_3_74),
       .pivot_in   (pivot_in_3_74),
       .start_out  (start_out_3_74),
       .swap_out   (swap_out_3_74),
       .data_out   (data_out_3_74),
       .op_out     (op_out_3_74),
       .pivot_out  (pivot_out_3_74),
       .r          (r_3_74)
     );

  // row 3, col 75

     reg start_in_3_75;
     wire start_out_3_75;

     reg swap_in_3_75;
     wire swap_out_3_75;

     reg [1:0] op_in_3_75;
     wire [1:0] op_out_3_75;

     wire r_3_75;

     reg data_in_3_75;
     wire data_out_3_75;

     reg pivot_in_3_75;
     wire pivot_out_3_75;

     always @(posedge clk) begin
         op_in_3_75 <= op_out_3_74;
         pivot_in_3_75 <= pivot_out_3_74;
         start_in_3_75 <= start_out_3_74;
         swap_in_3_75 <= swap_out_3_74;
     end

     always @(posedge clk) begin
         data_in_3_75 <= data_out_2_75;
     end
  
     processor_AB AB_3_75 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_75),
       .start_in   (start_in_3_75),
       .swap_in   (swap_in_3_75),
       .op_in      (op_in_3_75),
       .pivot_in   (pivot_in_3_75),
       .start_out  (start_out_3_75),
       .swap_out   (swap_out_3_75),
       .data_out   (data_out_3_75),
       .op_out     (op_out_3_75),
       .pivot_out  (pivot_out_3_75),
       .r          (r_3_75)
     );

  // row 3, col 76

     reg start_in_3_76;
     wire start_out_3_76;

     reg swap_in_3_76;
     wire swap_out_3_76;

     reg [1:0] op_in_3_76;
     wire [1:0] op_out_3_76;

     wire r_3_76;

     reg data_in_3_76;
     wire data_out_3_76;

     reg pivot_in_3_76;
     wire pivot_out_3_76;

     always @(posedge clk) begin
         op_in_3_76 <= op_out_3_75;
         pivot_in_3_76 <= pivot_out_3_75;
         start_in_3_76 <= start_out_3_75;
         swap_in_3_76 <= swap_out_3_75;
     end

     always @(posedge clk) begin
         data_in_3_76 <= data_out_2_76;
     end
  
     processor_AB AB_3_76 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_76),
       .start_in   (start_in_3_76),
       .swap_in   (swap_in_3_76),
       .op_in      (op_in_3_76),
       .pivot_in   (pivot_in_3_76),
       .start_out  (start_out_3_76),
       .swap_out   (swap_out_3_76),
       .data_out   (data_out_3_76),
       .op_out     (op_out_3_76),
       .pivot_out  (pivot_out_3_76),
       .r          (r_3_76)
     );

  // row 3, col 77

     reg start_in_3_77;
     wire start_out_3_77;

     reg swap_in_3_77;
     wire swap_out_3_77;

     reg [1:0] op_in_3_77;
     wire [1:0] op_out_3_77;

     wire r_3_77;

     reg data_in_3_77;
     wire data_out_3_77;

     reg pivot_in_3_77;
     wire pivot_out_3_77;

     always @(posedge clk) begin
         op_in_3_77 <= op_out_3_76;
         pivot_in_3_77 <= pivot_out_3_76;
         start_in_3_77 <= start_out_3_76;
         swap_in_3_77 <= swap_out_3_76;
     end

     always @(posedge clk) begin
         data_in_3_77 <= data_out_2_77;
     end
  
     processor_AB AB_3_77 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_77),
       .start_in   (start_in_3_77),
       .swap_in   (swap_in_3_77),
       .op_in      (op_in_3_77),
       .pivot_in   (pivot_in_3_77),
       .start_out  (start_out_3_77),
       .swap_out   (swap_out_3_77),
       .data_out   (data_out_3_77),
       .op_out     (op_out_3_77),
       .pivot_out  (pivot_out_3_77),
       .r          (r_3_77)
     );

  // row 3, col 78

     reg start_in_3_78;
     wire start_out_3_78;

     reg swap_in_3_78;
     wire swap_out_3_78;

     reg [1:0] op_in_3_78;
     wire [1:0] op_out_3_78;

     wire r_3_78;

     reg data_in_3_78;
     wire data_out_3_78;

     reg pivot_in_3_78;
     wire pivot_out_3_78;

     always @(posedge clk) begin
         op_in_3_78 <= op_out_3_77;
         pivot_in_3_78 <= pivot_out_3_77;
         start_in_3_78 <= start_out_3_77;
         swap_in_3_78 <= swap_out_3_77;
     end

     always @(posedge clk) begin
         data_in_3_78 <= data_out_2_78;
     end
  
     processor_AB AB_3_78 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_78),
       .start_in   (start_in_3_78),
       .swap_in   (swap_in_3_78),
       .op_in      (op_in_3_78),
       .pivot_in   (pivot_in_3_78),
       .start_out  (start_out_3_78),
       .swap_out   (swap_out_3_78),
       .data_out   (data_out_3_78),
       .op_out     (op_out_3_78),
       .pivot_out  (pivot_out_3_78),
       .r          (r_3_78)
     );

  // row 3, col 79

     reg start_in_3_79;
     wire start_out_3_79;

     reg swap_in_3_79;
     wire swap_out_3_79;

     reg [1:0] op_in_3_79;
     wire [1:0] op_out_3_79;

     wire r_3_79;

     reg data_in_3_79;
     wire data_out_3_79;

     reg pivot_in_3_79;
     wire pivot_out_3_79;

     always @(posedge clk) begin
         op_in_3_79 <= op_out_3_78;
         pivot_in_3_79 <= pivot_out_3_78;
         start_in_3_79 <= start_out_3_78;
         swap_in_3_79 <= swap_out_3_78;
     end

     always @(posedge clk) begin
         data_in_3_79 <= data_out_2_79;
     end
  
     processor_AB AB_3_79 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_79),
       .start_in   (start_in_3_79),
       .swap_in   (swap_in_3_79),
       .op_in      (op_in_3_79),
       .pivot_in   (pivot_in_3_79),
       .start_out  (start_out_3_79),
       .swap_out   (swap_out_3_79),
       .data_out   (data_out_3_79),
       .op_out     (op_out_3_79),
       .pivot_out  (pivot_out_3_79),
       .r          (r_3_79)
     );

  // row 3, col 80

     reg start_in_3_80;
     wire start_out_3_80;

     reg swap_in_3_80;
     wire swap_out_3_80;

     reg [1:0] op_in_3_80;
     wire [1:0] op_out_3_80;

     wire r_3_80;

     reg data_in_3_80;
     wire data_out_3_80;

     reg pivot_in_3_80;
     wire pivot_out_3_80;

     always @(posedge clk) begin
         op_in_3_80 <= op_out_3_79;
         pivot_in_3_80 <= pivot_out_3_79;
         start_in_3_80 <= start_out_3_79;
         swap_in_3_80 <= swap_out_3_79;
     end

     always @(posedge clk) begin
         data_in_3_80 <= data_out_2_80;
     end
  
     processor_AB AB_3_80 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_80),
       .start_in   (start_in_3_80),
       .swap_in   (swap_in_3_80),
       .op_in      (op_in_3_80),
       .pivot_in   (pivot_in_3_80),
       .start_out  (start_out_3_80),
       .swap_out   (swap_out_3_80),
       .data_out   (data_out_3_80),
       .op_out     (op_out_3_80),
       .pivot_out  (pivot_out_3_80),
       .r          (r_3_80)
     );

  // row 3, col 81

     reg start_in_3_81;
     wire start_out_3_81;

     reg swap_in_3_81;
     wire swap_out_3_81;

     reg [1:0] op_in_3_81;
     wire [1:0] op_out_3_81;

     wire r_3_81;

     reg data_in_3_81;
     wire data_out_3_81;

     reg pivot_in_3_81;
     wire pivot_out_3_81;

     always @(posedge clk) begin
         op_in_3_81 <= op_out_3_80;
         pivot_in_3_81 <= pivot_out_3_80;
         start_in_3_81 <= start_out_3_80;
         swap_in_3_81 <= swap_out_3_80;
     end

     always @(posedge clk) begin
         data_in_3_81 <= data_out_2_81;
     end
  
     processor_AB AB_3_81 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_81),
       .start_in   (start_in_3_81),
       .swap_in   (swap_in_3_81),
       .op_in      (op_in_3_81),
       .pivot_in   (pivot_in_3_81),
       .start_out  (start_out_3_81),
       .swap_out   (swap_out_3_81),
       .data_out   (data_out_3_81),
       .op_out     (op_out_3_81),
       .pivot_out  (pivot_out_3_81),
       .r          (r_3_81)
     );

  // row 3, col 82

     reg start_in_3_82;
     wire start_out_3_82;

     reg swap_in_3_82;
     wire swap_out_3_82;

     reg [1:0] op_in_3_82;
     wire [1:0] op_out_3_82;

     wire r_3_82;

     reg data_in_3_82;
     wire data_out_3_82;

     reg pivot_in_3_82;
     wire pivot_out_3_82;

     always @(posedge clk) begin
         op_in_3_82 <= op_out_3_81;
         pivot_in_3_82 <= pivot_out_3_81;
         start_in_3_82 <= start_out_3_81;
         swap_in_3_82 <= swap_out_3_81;
     end

     always @(posedge clk) begin
         data_in_3_82 <= data_out_2_82;
     end
  
     processor_AB AB_3_82 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_82),
       .start_in   (start_in_3_82),
       .swap_in   (swap_in_3_82),
       .op_in      (op_in_3_82),
       .pivot_in   (pivot_in_3_82),
       .start_out  (start_out_3_82),
       .swap_out   (swap_out_3_82),
       .data_out   (data_out_3_82),
       .op_out     (op_out_3_82),
       .pivot_out  (pivot_out_3_82),
       .r          (r_3_82)
     );

  // row 3, col 83

     reg start_in_3_83;
     wire start_out_3_83;

     reg swap_in_3_83;
     wire swap_out_3_83;

     reg [1:0] op_in_3_83;
     wire [1:0] op_out_3_83;

     wire r_3_83;

     reg data_in_3_83;
     wire data_out_3_83;

     reg pivot_in_3_83;
     wire pivot_out_3_83;

     always @(posedge clk) begin
         op_in_3_83 <= op_out_3_82;
         pivot_in_3_83 <= pivot_out_3_82;
         start_in_3_83 <= start_out_3_82;
         swap_in_3_83 <= swap_out_3_82;
     end

     always @(posedge clk) begin
         data_in_3_83 <= data_out_2_83;
     end
  
     processor_AB AB_3_83 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_83),
       .start_in   (start_in_3_83),
       .swap_in   (swap_in_3_83),
       .op_in      (op_in_3_83),
       .pivot_in   (pivot_in_3_83),
       .start_out  (start_out_3_83),
       .swap_out   (swap_out_3_83),
       .data_out   (data_out_3_83),
       .op_out     (op_out_3_83),
       .pivot_out  (pivot_out_3_83),
       .r          (r_3_83)
     );

  // row 3, col 84

     reg start_in_3_84;
     wire start_out_3_84;

     reg swap_in_3_84;
     wire swap_out_3_84;

     reg [1:0] op_in_3_84;
     wire [1:0] op_out_3_84;

     wire r_3_84;

     reg data_in_3_84;
     wire data_out_3_84;

     reg pivot_in_3_84;
     wire pivot_out_3_84;

     always @(posedge clk) begin
         op_in_3_84 <= op_out_3_83;
         pivot_in_3_84 <= pivot_out_3_83;
         start_in_3_84 <= start_out_3_83;
         swap_in_3_84 <= swap_out_3_83;
     end

     always @(posedge clk) begin
         data_in_3_84 <= data_out_2_84;
     end
  
     processor_AB AB_3_84 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_84),
       .start_in   (start_in_3_84),
       .swap_in   (swap_in_3_84),
       .op_in      (op_in_3_84),
       .pivot_in   (pivot_in_3_84),
       .start_out  (start_out_3_84),
       .swap_out   (swap_out_3_84),
       .data_out   (data_out_3_84),
       .op_out     (op_out_3_84),
       .pivot_out  (pivot_out_3_84),
       .r          (r_3_84)
     );

  // row 3, col 85

     reg start_in_3_85;
     wire start_out_3_85;

     reg swap_in_3_85;
     wire swap_out_3_85;

     reg [1:0] op_in_3_85;
     wire [1:0] op_out_3_85;

     wire r_3_85;

     reg data_in_3_85;
     wire data_out_3_85;

     reg pivot_in_3_85;
     wire pivot_out_3_85;

     always @(posedge clk) begin
         op_in_3_85 <= op_out_3_84;
         pivot_in_3_85 <= pivot_out_3_84;
         start_in_3_85 <= start_out_3_84;
         swap_in_3_85 <= swap_out_3_84;
     end

     always @(posedge clk) begin
         data_in_3_85 <= data_out_2_85;
     end
  
     processor_AB AB_3_85 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_85),
       .start_in   (start_in_3_85),
       .swap_in   (swap_in_3_85),
       .op_in      (op_in_3_85),
       .pivot_in   (pivot_in_3_85),
       .start_out  (start_out_3_85),
       .swap_out   (swap_out_3_85),
       .data_out   (data_out_3_85),
       .op_out     (op_out_3_85),
       .pivot_out  (pivot_out_3_85),
       .r          (r_3_85)
     );

  // row 3, col 86

     reg start_in_3_86;
     wire start_out_3_86;

     reg swap_in_3_86;
     wire swap_out_3_86;

     reg [1:0] op_in_3_86;
     wire [1:0] op_out_3_86;

     wire r_3_86;

     reg data_in_3_86;
     wire data_out_3_86;

     reg pivot_in_3_86;
     wire pivot_out_3_86;

     always @(posedge clk) begin
         op_in_3_86 <= op_out_3_85;
         pivot_in_3_86 <= pivot_out_3_85;
         start_in_3_86 <= start_out_3_85;
         swap_in_3_86 <= swap_out_3_85;
     end

     always @(posedge clk) begin
         data_in_3_86 <= data_out_2_86;
     end
  
     processor_AB AB_3_86 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_86),
       .start_in   (start_in_3_86),
       .swap_in   (swap_in_3_86),
       .op_in      (op_in_3_86),
       .pivot_in   (pivot_in_3_86),
       .start_out  (start_out_3_86),
       .swap_out   (swap_out_3_86),
       .data_out   (data_out_3_86),
       .op_out     (op_out_3_86),
       .pivot_out  (pivot_out_3_86),
       .r          (r_3_86)
     );

  // row 3, col 87

     reg start_in_3_87;
     wire start_out_3_87;

     reg swap_in_3_87;
     wire swap_out_3_87;

     reg [1:0] op_in_3_87;
     wire [1:0] op_out_3_87;

     wire r_3_87;

     reg data_in_3_87;
     wire data_out_3_87;

     reg pivot_in_3_87;
     wire pivot_out_3_87;

     always @(posedge clk) begin
         op_in_3_87 <= op_out_3_86;
         pivot_in_3_87 <= pivot_out_3_86;
         start_in_3_87 <= start_out_3_86;
         swap_in_3_87 <= swap_out_3_86;
     end

     always @(posedge clk) begin
         data_in_3_87 <= data_out_2_87;
     end
  
     processor_AB AB_3_87 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_87),
       .start_in   (start_in_3_87),
       .swap_in   (swap_in_3_87),
       .op_in      (op_in_3_87),
       .pivot_in   (pivot_in_3_87),
       .start_out  (start_out_3_87),
       .swap_out   (swap_out_3_87),
       .data_out   (data_out_3_87),
       .op_out     (op_out_3_87),
       .pivot_out  (pivot_out_3_87),
       .r          (r_3_87)
     );

  // row 3, col 88

     reg start_in_3_88;
     wire start_out_3_88;

     reg swap_in_3_88;
     wire swap_out_3_88;

     reg [1:0] op_in_3_88;
     wire [1:0] op_out_3_88;

     wire r_3_88;

     reg data_in_3_88;
     wire data_out_3_88;

     reg pivot_in_3_88;
     wire pivot_out_3_88;

     always @(posedge clk) begin
         op_in_3_88 <= op_out_3_87;
         pivot_in_3_88 <= pivot_out_3_87;
         start_in_3_88 <= start_out_3_87;
         swap_in_3_88 <= swap_out_3_87;
     end

     always @(posedge clk) begin
         data_in_3_88 <= data_out_2_88;
     end
  
     processor_AB AB_3_88 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_88),
       .start_in   (start_in_3_88),
       .swap_in   (swap_in_3_88),
       .op_in      (op_in_3_88),
       .pivot_in   (pivot_in_3_88),
       .start_out  (start_out_3_88),
       .swap_out   (swap_out_3_88),
       .data_out   (data_out_3_88),
       .op_out     (op_out_3_88),
       .pivot_out  (pivot_out_3_88),
       .r          (r_3_88)
     );

  // row 3, col 89

     reg start_in_3_89;
     wire start_out_3_89;

     reg swap_in_3_89;
     wire swap_out_3_89;

     reg [1:0] op_in_3_89;
     wire [1:0] op_out_3_89;

     wire r_3_89;

     reg data_in_3_89;
     wire data_out_3_89;

     reg pivot_in_3_89;
     wire pivot_out_3_89;

     always @(posedge clk) begin
         op_in_3_89 <= op_out_3_88;
         pivot_in_3_89 <= pivot_out_3_88;
         start_in_3_89 <= start_out_3_88;
         swap_in_3_89 <= swap_out_3_88;
     end

     always @(posedge clk) begin
         data_in_3_89 <= data_out_2_89;
     end
  
     processor_AB AB_3_89 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_89),
       .start_in   (start_in_3_89),
       .swap_in   (swap_in_3_89),
       .op_in      (op_in_3_89),
       .pivot_in   (pivot_in_3_89),
       .start_out  (start_out_3_89),
       .swap_out   (swap_out_3_89),
       .data_out   (data_out_3_89),
       .op_out     (op_out_3_89),
       .pivot_out  (pivot_out_3_89),
       .r          (r_3_89)
     );

  // row 3, col 90

     reg start_in_3_90;
     wire start_out_3_90;

     reg swap_in_3_90;
     wire swap_out_3_90;

     reg [1:0] op_in_3_90;
     wire [1:0] op_out_3_90;

     wire r_3_90;

     reg data_in_3_90;
     wire data_out_3_90;

     reg pivot_in_3_90;
     wire pivot_out_3_90;

     always @(posedge clk) begin
         op_in_3_90 <= op_out_3_89;
         pivot_in_3_90 <= pivot_out_3_89;
         start_in_3_90 <= start_out_3_89;
         swap_in_3_90 <= swap_out_3_89;
     end

     always @(posedge clk) begin
         data_in_3_90 <= data_out_2_90;
     end
  
     processor_AB AB_3_90 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_90),
       .start_in   (start_in_3_90),
       .swap_in   (swap_in_3_90),
       .op_in      (op_in_3_90),
       .pivot_in   (pivot_in_3_90),
       .start_out  (start_out_3_90),
       .swap_out   (swap_out_3_90),
       .data_out   (data_out_3_90),
       .op_out     (op_out_3_90),
       .pivot_out  (pivot_out_3_90),
       .r          (r_3_90)
     );

  // row 3, col 91

     reg start_in_3_91;
     wire start_out_3_91;

     reg swap_in_3_91;
     wire swap_out_3_91;

     reg [1:0] op_in_3_91;
     wire [1:0] op_out_3_91;

     wire r_3_91;

     reg data_in_3_91;
     wire data_out_3_91;

     reg pivot_in_3_91;
     wire pivot_out_3_91;

     always @(posedge clk) begin
         op_in_3_91 <= op_out_3_90;
         pivot_in_3_91 <= pivot_out_3_90;
         start_in_3_91 <= start_out_3_90;
         swap_in_3_91 <= swap_out_3_90;
     end

     always @(posedge clk) begin
         data_in_3_91 <= data_out_2_91;
     end
  
     processor_AB AB_3_91 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_91),
       .start_in   (start_in_3_91),
       .swap_in   (swap_in_3_91),
       .op_in      (op_in_3_91),
       .pivot_in   (pivot_in_3_91),
       .start_out  (start_out_3_91),
       .swap_out   (swap_out_3_91),
       .data_out   (data_out_3_91),
       .op_out     (op_out_3_91),
       .pivot_out  (pivot_out_3_91),
       .r          (r_3_91)
     );

  // row 3, col 92

     reg start_in_3_92;
     wire start_out_3_92;

     reg swap_in_3_92;
     wire swap_out_3_92;

     reg [1:0] op_in_3_92;
     wire [1:0] op_out_3_92;

     wire r_3_92;

     reg data_in_3_92;
     wire data_out_3_92;

     reg pivot_in_3_92;
     wire pivot_out_3_92;

     always @(posedge clk) begin
         op_in_3_92 <= op_out_3_91;
         pivot_in_3_92 <= pivot_out_3_91;
         start_in_3_92 <= start_out_3_91;
         swap_in_3_92 <= swap_out_3_91;
     end

     always @(posedge clk) begin
         data_in_3_92 <= data_out_2_92;
     end
  
     processor_AB AB_3_92 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_92),
       .start_in   (start_in_3_92),
       .swap_in   (swap_in_3_92),
       .op_in      (op_in_3_92),
       .pivot_in   (pivot_in_3_92),
       .start_out  (start_out_3_92),
       .swap_out   (swap_out_3_92),
       .data_out   (data_out_3_92),
       .op_out     (op_out_3_92),
       .pivot_out  (pivot_out_3_92),
       .r          (r_3_92)
     );

  // row 3, col 93

     reg start_in_3_93;
     wire start_out_3_93;

     reg swap_in_3_93;
     wire swap_out_3_93;

     reg [1:0] op_in_3_93;
     wire [1:0] op_out_3_93;

     wire r_3_93;

     reg data_in_3_93;
     wire data_out_3_93;

     reg pivot_in_3_93;
     wire pivot_out_3_93;

     always @(posedge clk) begin
         op_in_3_93 <= op_out_3_92;
         pivot_in_3_93 <= pivot_out_3_92;
         start_in_3_93 <= start_out_3_92;
         swap_in_3_93 <= swap_out_3_92;
     end

     always @(posedge clk) begin
         data_in_3_93 <= data_out_2_93;
     end
  
     processor_AB AB_3_93 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_93),
       .start_in   (start_in_3_93),
       .swap_in   (swap_in_3_93),
       .op_in      (op_in_3_93),
       .pivot_in   (pivot_in_3_93),
       .start_out  (start_out_3_93),
       .swap_out   (swap_out_3_93),
       .data_out   (data_out_3_93),
       .op_out     (op_out_3_93),
       .pivot_out  (pivot_out_3_93),
       .r          (r_3_93)
     );

  // row 3, col 94

     reg start_in_3_94;
     wire start_out_3_94;

     reg swap_in_3_94;
     wire swap_out_3_94;

     reg [1:0] op_in_3_94;
     wire [1:0] op_out_3_94;

     wire r_3_94;

     reg data_in_3_94;
     wire data_out_3_94;

     reg pivot_in_3_94;
     wire pivot_out_3_94;

     always @(posedge clk) begin
         op_in_3_94 <= op_out_3_93;
         pivot_in_3_94 <= pivot_out_3_93;
         start_in_3_94 <= start_out_3_93;
         swap_in_3_94 <= swap_out_3_93;
     end

     always @(posedge clk) begin
         data_in_3_94 <= data_out_2_94;
     end
  
     processor_AB AB_3_94 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_94),
       .start_in   (start_in_3_94),
       .swap_in   (swap_in_3_94),
       .op_in      (op_in_3_94),
       .pivot_in   (pivot_in_3_94),
       .start_out  (start_out_3_94),
       .swap_out   (swap_out_3_94),
       .data_out   (data_out_3_94),
       .op_out     (op_out_3_94),
       .pivot_out  (pivot_out_3_94),
       .r          (r_3_94)
     );

  // row 3, col 95

     reg start_in_3_95;
     wire start_out_3_95;

     reg swap_in_3_95;
     wire swap_out_3_95;

     reg [1:0] op_in_3_95;
     wire [1:0] op_out_3_95;

     wire r_3_95;

     reg data_in_3_95;
     wire data_out_3_95;

     reg pivot_in_3_95;
     wire pivot_out_3_95;

     always @(posedge clk) begin
         op_in_3_95 <= op_out_3_94;
         pivot_in_3_95 <= pivot_out_3_94;
         start_in_3_95 <= start_out_3_94;
         swap_in_3_95 <= swap_out_3_94;
     end

     always @(posedge clk) begin
         data_in_3_95 <= data_out_2_95;
     end
  
     processor_AB AB_3_95 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_95),
       .start_in   (start_in_3_95),
       .swap_in   (swap_in_3_95),
       .op_in      (op_in_3_95),
       .pivot_in   (pivot_in_3_95),
       .start_out  (start_out_3_95),
       .swap_out   (swap_out_3_95),
       .data_out   (data_out_3_95),
       .op_out     (op_out_3_95),
       .pivot_out  (pivot_out_3_95),
       .r          (r_3_95)
     );

  // row 3, col 96

     reg start_in_3_96;
     wire start_out_3_96;

     reg swap_in_3_96;
     wire swap_out_3_96;

     reg [1:0] op_in_3_96;
     wire [1:0] op_out_3_96;

     wire r_3_96;

     reg data_in_3_96;
     wire data_out_3_96;

     reg pivot_in_3_96;
     wire pivot_out_3_96;

     always @(posedge clk) begin
         op_in_3_96 <= op_out_3_95;
         pivot_in_3_96 <= pivot_out_3_95;
         start_in_3_96 <= start_out_3_95;
         swap_in_3_96 <= swap_out_3_95;
     end

     always @(posedge clk) begin
         data_in_3_96 <= data_out_2_96;
     end
  
     processor_AB AB_3_96 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_96),
       .start_in   (start_in_3_96),
       .swap_in   (swap_in_3_96),
       .op_in      (op_in_3_96),
       .pivot_in   (pivot_in_3_96),
       .start_out  (start_out_3_96),
       .swap_out   (swap_out_3_96),
       .data_out   (data_out_3_96),
       .op_out     (op_out_3_96),
       .pivot_out  (pivot_out_3_96),
       .r          (r_3_96)
     );

  // row 3, col 97

     reg start_in_3_97;
     wire start_out_3_97;

     reg swap_in_3_97;
     wire swap_out_3_97;

     reg [1:0] op_in_3_97;
     wire [1:0] op_out_3_97;

     wire r_3_97;

     reg data_in_3_97;
     wire data_out_3_97;

     reg pivot_in_3_97;
     wire pivot_out_3_97;

     always @(posedge clk) begin
         op_in_3_97 <= op_out_3_96;
         pivot_in_3_97 <= pivot_out_3_96;
         start_in_3_97 <= start_out_3_96;
         swap_in_3_97 <= swap_out_3_96;
     end

     always @(posedge clk) begin
         data_in_3_97 <= data_out_2_97;
     end
  
     processor_AB AB_3_97 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_97),
       .start_in   (start_in_3_97),
       .swap_in   (swap_in_3_97),
       .op_in      (op_in_3_97),
       .pivot_in   (pivot_in_3_97),
       .start_out  (start_out_3_97),
       .swap_out   (swap_out_3_97),
       .data_out   (data_out_3_97),
       .op_out     (op_out_3_97),
       .pivot_out  (pivot_out_3_97),
       .r          (r_3_97)
     );

  // row 3, col 98

     reg start_in_3_98;
     wire start_out_3_98;

     reg swap_in_3_98;
     wire swap_out_3_98;

     reg [1:0] op_in_3_98;
     wire [1:0] op_out_3_98;

     wire r_3_98;

     reg data_in_3_98;
     wire data_out_3_98;

     reg pivot_in_3_98;
     wire pivot_out_3_98;

     always @(posedge clk) begin
         op_in_3_98 <= op_out_3_97;
         pivot_in_3_98 <= pivot_out_3_97;
         start_in_3_98 <= start_out_3_97;
         swap_in_3_98 <= swap_out_3_97;
     end

     always @(posedge clk) begin
         data_in_3_98 <= data_out_2_98;
     end
  
     processor_AB AB_3_98 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_98),
       .start_in   (start_in_3_98),
       .swap_in   (swap_in_3_98),
       .op_in      (op_in_3_98),
       .pivot_in   (pivot_in_3_98),
       .start_out  (start_out_3_98),
       .swap_out   (swap_out_3_98),
       .data_out   (data_out_3_98),
       .op_out     (op_out_3_98),
       .pivot_out  (pivot_out_3_98),
       .r          (r_3_98)
     );

  // row 3, col 99

     reg start_in_3_99;
     wire start_out_3_99;

     reg swap_in_3_99;
     wire swap_out_3_99;

     reg [1:0] op_in_3_99;
     wire [1:0] op_out_3_99;

     wire r_3_99;

     reg data_in_3_99;
     wire data_out_3_99;

     reg pivot_in_3_99;
     wire pivot_out_3_99;

     always @(posedge clk) begin
         op_in_3_99 <= op_out_3_98;
         pivot_in_3_99 <= pivot_out_3_98;
         start_in_3_99 <= start_out_3_98;
         swap_in_3_99 <= swap_out_3_98;
     end

     always @(posedge clk) begin
         data_in_3_99 <= data_out_2_99;
     end
  
     processor_AB AB_3_99 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_99),
       .start_in   (start_in_3_99),
       .swap_in   (swap_in_3_99),
       .op_in      (op_in_3_99),
       .pivot_in   (pivot_in_3_99),
       .start_out  (start_out_3_99),
       .swap_out   (swap_out_3_99),
       .data_out   (data_out_3_99),
       .op_out     (op_out_3_99),
       .pivot_out  (pivot_out_3_99),
       .r          (r_3_99)
     );

  // row 3, col 100

     reg start_in_3_100;
     wire start_out_3_100;

     reg swap_in_3_100;
     wire swap_out_3_100;

     reg [1:0] op_in_3_100;
     wire [1:0] op_out_3_100;

     wire r_3_100;

     reg data_in_3_100;
     wire data_out_3_100;

     reg pivot_in_3_100;
     wire pivot_out_3_100;

     always @(posedge clk) begin
         op_in_3_100 <= op_out_3_99;
         pivot_in_3_100 <= pivot_out_3_99;
         start_in_3_100 <= start_out_3_99;
         swap_in_3_100 <= swap_out_3_99;
     end

     always @(posedge clk) begin
         data_in_3_100 <= data_out_2_100;
     end
  
     processor_AB AB_3_100 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_100),
       .start_in   (start_in_3_100),
       .swap_in   (swap_in_3_100),
       .op_in      (op_in_3_100),
       .pivot_in   (pivot_in_3_100),
       .start_out  (start_out_3_100),
       .swap_out   (swap_out_3_100),
       .data_out   (data_out_3_100),
       .op_out     (op_out_3_100),
       .pivot_out  (pivot_out_3_100),
       .r          (r_3_100)
     );

  // row 3, col 101

     reg start_in_3_101;
     wire start_out_3_101;

     reg swap_in_3_101;
     wire swap_out_3_101;

     reg [1:0] op_in_3_101;
     wire [1:0] op_out_3_101;

     wire r_3_101;

     reg data_in_3_101;
     wire data_out_3_101;

     reg pivot_in_3_101;
     wire pivot_out_3_101;

     always @(posedge clk) begin
         op_in_3_101 <= op_out_3_100;
         pivot_in_3_101 <= pivot_out_3_100;
         start_in_3_101 <= start_out_3_100;
         swap_in_3_101 <= swap_out_3_100;
     end

     always @(posedge clk) begin
         data_in_3_101 <= data_out_2_101;
     end
  
     processor_AB AB_3_101 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_101),
       .start_in   (start_in_3_101),
       .swap_in   (swap_in_3_101),
       .op_in      (op_in_3_101),
       .pivot_in   (pivot_in_3_101),
       .start_out  (start_out_3_101),
       .swap_out   (swap_out_3_101),
       .data_out   (data_out_3_101),
       .op_out     (op_out_3_101),
       .pivot_out  (pivot_out_3_101),
       .r          (r_3_101)
     );

  // row 3, col 102

     reg start_in_3_102;
     wire start_out_3_102;

     reg swap_in_3_102;
     wire swap_out_3_102;

     reg [1:0] op_in_3_102;
     wire [1:0] op_out_3_102;

     wire r_3_102;

     reg data_in_3_102;
     wire data_out_3_102;

     reg pivot_in_3_102;
     wire pivot_out_3_102;

     always @(posedge clk) begin
         op_in_3_102 <= op_out_3_101;
         pivot_in_3_102 <= pivot_out_3_101;
         start_in_3_102 <= start_out_3_101;
         swap_in_3_102 <= swap_out_3_101;
     end

     always @(posedge clk) begin
         data_in_3_102 <= data_out_2_102;
     end
  
     processor_AB AB_3_102 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_102),
       .start_in   (start_in_3_102),
       .swap_in   (swap_in_3_102),
       .op_in      (op_in_3_102),
       .pivot_in   (pivot_in_3_102),
       .start_out  (start_out_3_102),
       .swap_out   (swap_out_3_102),
       .data_out   (data_out_3_102),
       .op_out     (op_out_3_102),
       .pivot_out  (pivot_out_3_102),
       .r          (r_3_102)
     );

  // row 3, col 103

     reg start_in_3_103;
     wire start_out_3_103;

     reg swap_in_3_103;
     wire swap_out_3_103;

     reg [1:0] op_in_3_103;
     wire [1:0] op_out_3_103;

     wire r_3_103;

     reg data_in_3_103;
     wire data_out_3_103;

     reg pivot_in_3_103;
     wire pivot_out_3_103;

     always @(posedge clk) begin
         op_in_3_103 <= op_out_3_102;
         pivot_in_3_103 <= pivot_out_3_102;
         start_in_3_103 <= start_out_3_102;
         swap_in_3_103 <= swap_out_3_102;
     end

     always @(posedge clk) begin
         data_in_3_103 <= data_out_2_103;
     end
  
     processor_AB AB_3_103 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_103),
       .start_in   (start_in_3_103),
       .swap_in   (swap_in_3_103),
       .op_in      (op_in_3_103),
       .pivot_in   (pivot_in_3_103),
       .start_out  (start_out_3_103),
       .swap_out   (swap_out_3_103),
       .data_out   (data_out_3_103),
       .op_out     (op_out_3_103),
       .pivot_out  (pivot_out_3_103),
       .r          (r_3_103)
     );

  // row 3, col 104

     reg start_in_3_104;
     wire start_out_3_104;

     reg swap_in_3_104;
     wire swap_out_3_104;

     reg [1:0] op_in_3_104;
     wire [1:0] op_out_3_104;

     wire r_3_104;

     reg data_in_3_104;
     wire data_out_3_104;

     reg pivot_in_3_104;
     wire pivot_out_3_104;

     always @(posedge clk) begin
         op_in_3_104 <= op_out_3_103;
         pivot_in_3_104 <= pivot_out_3_103;
         start_in_3_104 <= start_out_3_103;
         swap_in_3_104 <= swap_out_3_103;
     end

     always @(posedge clk) begin
         data_in_3_104 <= data_out_2_104;
     end
  
     processor_AB AB_3_104 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_104),
       .start_in   (start_in_3_104),
       .swap_in   (swap_in_3_104),
       .op_in      (op_in_3_104),
       .pivot_in   (pivot_in_3_104),
       .start_out  (start_out_3_104),
       .swap_out   (swap_out_3_104),
       .data_out   (data_out_3_104),
       .op_out     (op_out_3_104),
       .pivot_out  (pivot_out_3_104),
       .r          (r_3_104)
     );

  // row 3, col 105

     reg start_in_3_105;
     wire start_out_3_105;

     reg swap_in_3_105;
     wire swap_out_3_105;

     reg [1:0] op_in_3_105;
     wire [1:0] op_out_3_105;

     wire r_3_105;

     reg data_in_3_105;
     wire data_out_3_105;

     reg pivot_in_3_105;
     wire pivot_out_3_105;

     always @(posedge clk) begin
         op_in_3_105 <= op_out_3_104;
         pivot_in_3_105 <= pivot_out_3_104;
         start_in_3_105 <= start_out_3_104;
         swap_in_3_105 <= swap_out_3_104;
     end

     always @(posedge clk) begin
         data_in_3_105 <= data_out_2_105;
     end
  
     processor_AB AB_3_105 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_105),
       .start_in   (start_in_3_105),
       .swap_in   (swap_in_3_105),
       .op_in      (op_in_3_105),
       .pivot_in   (pivot_in_3_105),
       .start_out  (start_out_3_105),
       .swap_out   (swap_out_3_105),
       .data_out   (data_out_3_105),
       .op_out     (op_out_3_105),
       .pivot_out  (pivot_out_3_105),
       .r          (r_3_105)
     );

  // row 3, col 106

     reg start_in_3_106;
     wire start_out_3_106;

     reg swap_in_3_106;
     wire swap_out_3_106;

     reg [1:0] op_in_3_106;
     wire [1:0] op_out_3_106;

     wire r_3_106;

     reg data_in_3_106;
     wire data_out_3_106;

     reg pivot_in_3_106;
     wire pivot_out_3_106;

     always @(posedge clk) begin
         op_in_3_106 <= op_out_3_105;
         pivot_in_3_106 <= pivot_out_3_105;
         start_in_3_106 <= start_out_3_105;
         swap_in_3_106 <= swap_out_3_105;
     end

     always @(posedge clk) begin
         data_in_3_106 <= data_out_2_106;
     end
  
     processor_AB AB_3_106 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_106),
       .start_in   (start_in_3_106),
       .swap_in   (swap_in_3_106),
       .op_in      (op_in_3_106),
       .pivot_in   (pivot_in_3_106),
       .start_out  (start_out_3_106),
       .swap_out   (swap_out_3_106),
       .data_out   (data_out_3_106),
       .op_out     (op_out_3_106),
       .pivot_out  (pivot_out_3_106),
       .r          (r_3_106)
     );

  // row 3, col 107

     reg start_in_3_107;
     wire start_out_3_107;

     reg swap_in_3_107;
     wire swap_out_3_107;

     reg [1:0] op_in_3_107;
     wire [1:0] op_out_3_107;

     wire r_3_107;

     reg data_in_3_107;
     wire data_out_3_107;

     reg pivot_in_3_107;
     wire pivot_out_3_107;

     always @(posedge clk) begin
         op_in_3_107 <= op_out_3_106;
         pivot_in_3_107 <= pivot_out_3_106;
         start_in_3_107 <= start_out_3_106;
         swap_in_3_107 <= swap_out_3_106;
     end

     always @(posedge clk) begin
         data_in_3_107 <= data_out_2_107;
     end
  
     processor_AB AB_3_107 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_107),
       .start_in   (start_in_3_107),
       .swap_in   (swap_in_3_107),
       .op_in      (op_in_3_107),
       .pivot_in   (pivot_in_3_107),
       .start_out  (start_out_3_107),
       .swap_out   (swap_out_3_107),
       .data_out   (data_out_3_107),
       .op_out     (op_out_3_107),
       .pivot_out  (pivot_out_3_107),
       .r          (r_3_107)
     );

  // row 3, col 108

     reg start_in_3_108;
     wire start_out_3_108;

     reg swap_in_3_108;
     wire swap_out_3_108;

     reg [1:0] op_in_3_108;
     wire [1:0] op_out_3_108;

     wire r_3_108;

     reg data_in_3_108;
     wire data_out_3_108;

     reg pivot_in_3_108;
     wire pivot_out_3_108;

     always @(posedge clk) begin
         op_in_3_108 <= op_out_3_107;
         pivot_in_3_108 <= pivot_out_3_107;
         start_in_3_108 <= start_out_3_107;
         swap_in_3_108 <= swap_out_3_107;
     end

     always @(posedge clk) begin
         data_in_3_108 <= data_out_2_108;
     end
  
     processor_AB AB_3_108 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_108),
       .start_in   (start_in_3_108),
       .swap_in   (swap_in_3_108),
       .op_in      (op_in_3_108),
       .pivot_in   (pivot_in_3_108),
       .start_out  (start_out_3_108),
       .swap_out   (swap_out_3_108),
       .data_out   (data_out_3_108),
       .op_out     (op_out_3_108),
       .pivot_out  (pivot_out_3_108),
       .r          (r_3_108)
     );

  // row 3, col 109

     reg start_in_3_109;
     wire start_out_3_109;

     reg swap_in_3_109;
     wire swap_out_3_109;

     reg [1:0] op_in_3_109;
     wire [1:0] op_out_3_109;

     wire r_3_109;

     reg data_in_3_109;
     wire data_out_3_109;

     reg pivot_in_3_109;
     wire pivot_out_3_109;

     always @(posedge clk) begin
         op_in_3_109 <= op_out_3_108;
         pivot_in_3_109 <= pivot_out_3_108;
         start_in_3_109 <= start_out_3_108;
         swap_in_3_109 <= swap_out_3_108;
     end

     always @(posedge clk) begin
         data_in_3_109 <= data_out_2_109;
     end
  
     processor_AB AB_3_109 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_109),
       .start_in   (start_in_3_109),
       .swap_in   (swap_in_3_109),
       .op_in      (op_in_3_109),
       .pivot_in   (pivot_in_3_109),
       .start_out  (start_out_3_109),
       .swap_out   (swap_out_3_109),
       .data_out   (data_out_3_109),
       .op_out     (op_out_3_109),
       .pivot_out  (pivot_out_3_109),
       .r          (r_3_109)
     );

  // row 3, col 110

     reg start_in_3_110;
     wire start_out_3_110;

     reg swap_in_3_110;
     wire swap_out_3_110;

     reg [1:0] op_in_3_110;
     wire [1:0] op_out_3_110;

     wire r_3_110;

     reg data_in_3_110;
     wire data_out_3_110;

     reg pivot_in_3_110;
     wire pivot_out_3_110;

     always @(posedge clk) begin
         op_in_3_110 <= op_out_3_109;
         pivot_in_3_110 <= pivot_out_3_109;
         start_in_3_110 <= start_out_3_109;
         swap_in_3_110 <= swap_out_3_109;
     end

     always @(posedge clk) begin
         data_in_3_110 <= data_out_2_110;
     end
  
     processor_AB AB_3_110 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_110),
       .start_in   (start_in_3_110),
       .swap_in   (swap_in_3_110),
       .op_in      (op_in_3_110),
       .pivot_in   (pivot_in_3_110),
       .start_out  (start_out_3_110),
       .swap_out   (swap_out_3_110),
       .data_out   (data_out_3_110),
       .op_out     (op_out_3_110),
       .pivot_out  (pivot_out_3_110),
       .r          (r_3_110)
     );

  // row 3, col 111

     reg start_in_3_111;
     wire start_out_3_111;

     reg swap_in_3_111;
     wire swap_out_3_111;

     reg [1:0] op_in_3_111;
     wire [1:0] op_out_3_111;

     wire r_3_111;

     reg data_in_3_111;
     wire data_out_3_111;

     reg pivot_in_3_111;
     wire pivot_out_3_111;

     always @(posedge clk) begin
         op_in_3_111 <= op_out_3_110;
         pivot_in_3_111 <= pivot_out_3_110;
         start_in_3_111 <= start_out_3_110;
         swap_in_3_111 <= swap_out_3_110;
     end

     always @(posedge clk) begin
         data_in_3_111 <= data_out_2_111;
     end
  
     processor_AB AB_3_111 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_111),
       .start_in   (start_in_3_111),
       .swap_in   (swap_in_3_111),
       .op_in      (op_in_3_111),
       .pivot_in   (pivot_in_3_111),
       .start_out  (start_out_3_111),
       .swap_out   (swap_out_3_111),
       .data_out   (data_out_3_111),
       .op_out     (op_out_3_111),
       .pivot_out  (pivot_out_3_111),
       .r          (r_3_111)
     );

  // row 3, col 112

     reg start_in_3_112;
     wire start_out_3_112;

     reg swap_in_3_112;
     wire swap_out_3_112;

     reg [1:0] op_in_3_112;
     wire [1:0] op_out_3_112;

     wire r_3_112;

     reg data_in_3_112;
     wire data_out_3_112;

     reg pivot_in_3_112;
     wire pivot_out_3_112;

     always @(posedge clk) begin
         op_in_3_112 <= op_out_3_111;
         pivot_in_3_112 <= pivot_out_3_111;
         start_in_3_112 <= start_out_3_111;
         swap_in_3_112 <= swap_out_3_111;
     end

     always @(posedge clk) begin
         data_in_3_112 <= data_out_2_112;
     end
  
     processor_AB AB_3_112 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_112),
       .start_in   (start_in_3_112),
       .swap_in   (swap_in_3_112),
       .op_in      (op_in_3_112),
       .pivot_in   (pivot_in_3_112),
       .start_out  (start_out_3_112),
       .swap_out   (swap_out_3_112),
       .data_out   (data_out_3_112),
       .op_out     (op_out_3_112),
       .pivot_out  (pivot_out_3_112),
       .r          (r_3_112)
     );

  // row 3, col 113

     reg start_in_3_113;
     wire start_out_3_113;

     reg swap_in_3_113;
     wire swap_out_3_113;

     reg [1:0] op_in_3_113;
     wire [1:0] op_out_3_113;

     wire r_3_113;

     reg data_in_3_113;
     wire data_out_3_113;

     reg pivot_in_3_113;
     wire pivot_out_3_113;

     always @(posedge clk) begin
         op_in_3_113 <= op_out_3_112;
         pivot_in_3_113 <= pivot_out_3_112;
         start_in_3_113 <= start_out_3_112;
         swap_in_3_113 <= swap_out_3_112;
     end

     always @(posedge clk) begin
         data_in_3_113 <= data_out_2_113;
     end
  
     processor_AB AB_3_113 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_113),
       .start_in   (start_in_3_113),
       .swap_in   (swap_in_3_113),
       .op_in      (op_in_3_113),
       .pivot_in   (pivot_in_3_113),
       .start_out  (start_out_3_113),
       .swap_out   (swap_out_3_113),
       .data_out   (data_out_3_113),
       .op_out     (op_out_3_113),
       .pivot_out  (pivot_out_3_113),
       .r          (r_3_113)
     );

  // row 3, col 114

     reg start_in_3_114;
     wire start_out_3_114;

     reg swap_in_3_114;
     wire swap_out_3_114;

     reg [1:0] op_in_3_114;
     wire [1:0] op_out_3_114;

     wire r_3_114;

     reg data_in_3_114;
     wire data_out_3_114;

     reg pivot_in_3_114;
     wire pivot_out_3_114;

     always @(posedge clk) begin
         op_in_3_114 <= op_out_3_113;
         pivot_in_3_114 <= pivot_out_3_113;
         start_in_3_114 <= start_out_3_113;
         swap_in_3_114 <= swap_out_3_113;
     end

     always @(posedge clk) begin
         data_in_3_114 <= data_out_2_114;
     end
  
     processor_AB AB_3_114 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_114),
       .start_in   (start_in_3_114),
       .swap_in   (swap_in_3_114),
       .op_in      (op_in_3_114),
       .pivot_in   (pivot_in_3_114),
       .start_out  (start_out_3_114),
       .swap_out   (swap_out_3_114),
       .data_out   (data_out_3_114),
       .op_out     (op_out_3_114),
       .pivot_out  (pivot_out_3_114),
       .r          (r_3_114)
     );

  // row 3, col 115

     reg start_in_3_115;
     wire start_out_3_115;

     reg swap_in_3_115;
     wire swap_out_3_115;

     reg [1:0] op_in_3_115;
     wire [1:0] op_out_3_115;

     wire r_3_115;

     reg data_in_3_115;
     wire data_out_3_115;

     reg pivot_in_3_115;
     wire pivot_out_3_115;

     always @(posedge clk) begin
         op_in_3_115 <= op_out_3_114;
         pivot_in_3_115 <= pivot_out_3_114;
         start_in_3_115 <= start_out_3_114;
         swap_in_3_115 <= swap_out_3_114;
     end

     always @(posedge clk) begin
         data_in_3_115 <= data_out_2_115;
     end
  
     processor_AB AB_3_115 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_115),
       .start_in   (start_in_3_115),
       .swap_in   (swap_in_3_115),
       .op_in      (op_in_3_115),
       .pivot_in   (pivot_in_3_115),
       .start_out  (start_out_3_115),
       .swap_out   (swap_out_3_115),
       .data_out   (data_out_3_115),
       .op_out     (op_out_3_115),
       .pivot_out  (pivot_out_3_115),
       .r          (r_3_115)
     );

  // row 3, col 116

     reg start_in_3_116;
     wire start_out_3_116;

     reg swap_in_3_116;
     wire swap_out_3_116;

     reg [1:0] op_in_3_116;
     wire [1:0] op_out_3_116;

     wire r_3_116;

     reg data_in_3_116;
     wire data_out_3_116;

     reg pivot_in_3_116;
     wire pivot_out_3_116;

     always @(posedge clk) begin
         op_in_3_116 <= op_out_3_115;
         pivot_in_3_116 <= pivot_out_3_115;
         start_in_3_116 <= start_out_3_115;
         swap_in_3_116 <= swap_out_3_115;
     end

     always @(posedge clk) begin
         data_in_3_116 <= data_out_2_116;
     end
  
     processor_AB AB_3_116 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_116),
       .start_in   (start_in_3_116),
       .swap_in   (swap_in_3_116),
       .op_in      (op_in_3_116),
       .pivot_in   (pivot_in_3_116),
       .start_out  (start_out_3_116),
       .swap_out   (swap_out_3_116),
       .data_out   (data_out_3_116),
       .op_out     (op_out_3_116),
       .pivot_out  (pivot_out_3_116),
       .r          (r_3_116)
     );

  // row 3, col 117

     reg start_in_3_117;
     wire start_out_3_117;

     reg swap_in_3_117;
     wire swap_out_3_117;

     reg [1:0] op_in_3_117;
     wire [1:0] op_out_3_117;

     wire r_3_117;

     reg data_in_3_117;
     wire data_out_3_117;

     reg pivot_in_3_117;
     wire pivot_out_3_117;

     always @(posedge clk) begin
         op_in_3_117 <= op_out_3_116;
         pivot_in_3_117 <= pivot_out_3_116;
         start_in_3_117 <= start_out_3_116;
         swap_in_3_117 <= swap_out_3_116;
     end

     always @(posedge clk) begin
         data_in_3_117 <= data_out_2_117;
     end
  
     processor_AB AB_3_117 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_117),
       .start_in   (start_in_3_117),
       .swap_in   (swap_in_3_117),
       .op_in      (op_in_3_117),
       .pivot_in   (pivot_in_3_117),
       .start_out  (start_out_3_117),
       .swap_out   (swap_out_3_117),
       .data_out   (data_out_3_117),
       .op_out     (op_out_3_117),
       .pivot_out  (pivot_out_3_117),
       .r          (r_3_117)
     );

  // row 3, col 118

     reg start_in_3_118;
     wire start_out_3_118;

     reg swap_in_3_118;
     wire swap_out_3_118;

     reg [1:0] op_in_3_118;
     wire [1:0] op_out_3_118;

     wire r_3_118;

     reg data_in_3_118;
     wire data_out_3_118;

     reg pivot_in_3_118;
     wire pivot_out_3_118;

     always @(posedge clk) begin
         op_in_3_118 <= op_out_3_117;
         pivot_in_3_118 <= pivot_out_3_117;
         start_in_3_118 <= start_out_3_117;
         swap_in_3_118 <= swap_out_3_117;
     end

     always @(posedge clk) begin
         data_in_3_118 <= data_out_2_118;
     end
  
     processor_AB AB_3_118 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_118),
       .start_in   (start_in_3_118),
       .swap_in   (swap_in_3_118),
       .op_in      (op_in_3_118),
       .pivot_in   (pivot_in_3_118),
       .start_out  (start_out_3_118),
       .swap_out   (swap_out_3_118),
       .data_out   (data_out_3_118),
       .op_out     (op_out_3_118),
       .pivot_out  (pivot_out_3_118),
       .r          (r_3_118)
     );

  // row 3, col 119

     reg start_in_3_119;
     wire start_out_3_119;

     reg swap_in_3_119;
     wire swap_out_3_119;

     reg [1:0] op_in_3_119;
     wire [1:0] op_out_3_119;

     wire r_3_119;

     reg data_in_3_119;
     wire data_out_3_119;

     reg pivot_in_3_119;
     wire pivot_out_3_119;

     always @(posedge clk) begin
         op_in_3_119 <= op_out_3_118;
         pivot_in_3_119 <= pivot_out_3_118;
         start_in_3_119 <= start_out_3_118;
         swap_in_3_119 <= swap_out_3_118;
     end

     always @(posedge clk) begin
         data_in_3_119 <= data_out_2_119;
     end
  
     processor_AB AB_3_119 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_119),
       .start_in   (start_in_3_119),
       .swap_in   (swap_in_3_119),
       .op_in      (op_in_3_119),
       .pivot_in   (pivot_in_3_119),
       .start_out  (start_out_3_119),
       .swap_out   (swap_out_3_119),
       .data_out   (data_out_3_119),
       .op_out     (op_out_3_119),
       .pivot_out  (pivot_out_3_119),
       .r          (r_3_119)
     );

  // row 3, col 120

     reg start_in_3_120;
     wire start_out_3_120;

     reg swap_in_3_120;
     wire swap_out_3_120;

     reg [1:0] op_in_3_120;
     wire [1:0] op_out_3_120;

     wire r_3_120;

     reg data_in_3_120;
     wire data_out_3_120;

     reg pivot_in_3_120;
     wire pivot_out_3_120;

     always @(posedge clk) begin
         op_in_3_120 <= op_out_3_119;
         pivot_in_3_120 <= pivot_out_3_119;
         start_in_3_120 <= start_out_3_119;
         swap_in_3_120 <= swap_out_3_119;
     end

     always @(posedge clk) begin
         data_in_3_120 <= data_out_2_120;
     end
  
     processor_AB AB_3_120 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_120),
       .start_in   (start_in_3_120),
       .swap_in   (swap_in_3_120),
       .op_in      (op_in_3_120),
       .pivot_in   (pivot_in_3_120),
       .start_out  (start_out_3_120),
       .swap_out   (swap_out_3_120),
       .data_out   (data_out_3_120),
       .op_out     (op_out_3_120),
       .pivot_out  (pivot_out_3_120),
       .r          (r_3_120)
     );

  // row 3, col 121

     reg start_in_3_121;
     wire start_out_3_121;

     reg swap_in_3_121;
     wire swap_out_3_121;

     reg [1:0] op_in_3_121;
     wire [1:0] op_out_3_121;

     wire r_3_121;

     reg data_in_3_121;
     wire data_out_3_121;

     reg pivot_in_3_121;
     wire pivot_out_3_121;

     always @(posedge clk) begin
         op_in_3_121 <= op_out_3_120;
         pivot_in_3_121 <= pivot_out_3_120;
         start_in_3_121 <= start_out_3_120;
         swap_in_3_121 <= swap_out_3_120;
     end

     always @(posedge clk) begin
         data_in_3_121 <= data_out_2_121;
     end
  
     processor_AB AB_3_121 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_121),
       .start_in   (start_in_3_121),
       .swap_in   (swap_in_3_121),
       .op_in      (op_in_3_121),
       .pivot_in   (pivot_in_3_121),
       .start_out  (start_out_3_121),
       .swap_out   (swap_out_3_121),
       .data_out   (data_out_3_121),
       .op_out     (op_out_3_121),
       .pivot_out  (pivot_out_3_121),
       .r          (r_3_121)
     );

  // row 3, col 122

     reg start_in_3_122;
     wire start_out_3_122;

     reg swap_in_3_122;
     wire swap_out_3_122;

     reg [1:0] op_in_3_122;
     wire [1:0] op_out_3_122;

     wire r_3_122;

     reg data_in_3_122;
     wire data_out_3_122;

     reg pivot_in_3_122;
     wire pivot_out_3_122;

     always @(posedge clk) begin
         op_in_3_122 <= op_out_3_121;
         pivot_in_3_122 <= pivot_out_3_121;
         start_in_3_122 <= start_out_3_121;
         swap_in_3_122 <= swap_out_3_121;
     end

     always @(posedge clk) begin
         data_in_3_122 <= data_out_2_122;
     end
  
     processor_AB AB_3_122 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_122),
       .start_in   (start_in_3_122),
       .swap_in   (swap_in_3_122),
       .op_in      (op_in_3_122),
       .pivot_in   (pivot_in_3_122),
       .start_out  (start_out_3_122),
       .swap_out   (swap_out_3_122),
       .data_out   (data_out_3_122),
       .op_out     (op_out_3_122),
       .pivot_out  (pivot_out_3_122),
       .r          (r_3_122)
     );

  // row 3, col 123

     reg start_in_3_123;
     wire start_out_3_123;

     reg swap_in_3_123;
     wire swap_out_3_123;

     reg [1:0] op_in_3_123;
     wire [1:0] op_out_3_123;

     wire r_3_123;

     reg data_in_3_123;
     wire data_out_3_123;

     reg pivot_in_3_123;
     wire pivot_out_3_123;

     always @(posedge clk) begin
         op_in_3_123 <= op_out_3_122;
         pivot_in_3_123 <= pivot_out_3_122;
         start_in_3_123 <= start_out_3_122;
         swap_in_3_123 <= swap_out_3_122;
     end

     always @(posedge clk) begin
         data_in_3_123 <= data_out_2_123;
     end
  
     processor_AB AB_3_123 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_123),
       .start_in   (start_in_3_123),
       .swap_in   (swap_in_3_123),
       .op_in      (op_in_3_123),
       .pivot_in   (pivot_in_3_123),
       .start_out  (start_out_3_123),
       .swap_out   (swap_out_3_123),
       .data_out   (data_out_3_123),
       .op_out     (op_out_3_123),
       .pivot_out  (pivot_out_3_123),
       .r          (r_3_123)
     );

  // row 3, col 124

     reg start_in_3_124;
     wire start_out_3_124;

     reg swap_in_3_124;
     wire swap_out_3_124;

     reg [1:0] op_in_3_124;
     wire [1:0] op_out_3_124;

     wire r_3_124;

     reg data_in_3_124;
     wire data_out_3_124;

     reg pivot_in_3_124;
     wire pivot_out_3_124;

     always @(posedge clk) begin
         op_in_3_124 <= op_out_3_123;
         pivot_in_3_124 <= pivot_out_3_123;
         start_in_3_124 <= start_out_3_123;
         swap_in_3_124 <= swap_out_3_123;
     end

     always @(posedge clk) begin
         data_in_3_124 <= data_out_2_124;
     end
  
     processor_AB AB_3_124 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_124),
       .start_in   (start_in_3_124),
       .swap_in   (swap_in_3_124),
       .op_in      (op_in_3_124),
       .pivot_in   (pivot_in_3_124),
       .start_out  (start_out_3_124),
       .swap_out   (swap_out_3_124),
       .data_out   (data_out_3_124),
       .op_out     (op_out_3_124),
       .pivot_out  (pivot_out_3_124),
       .r          (r_3_124)
     );

  // row 3, col 125

     reg start_in_3_125;
     wire start_out_3_125;

     reg swap_in_3_125;
     wire swap_out_3_125;

     reg [1:0] op_in_3_125;
     wire [1:0] op_out_3_125;

     wire r_3_125;

     reg data_in_3_125;
     wire data_out_3_125;

     reg pivot_in_3_125;
     wire pivot_out_3_125;

     always @(posedge clk) begin
         op_in_3_125 <= op_out_3_124;
         pivot_in_3_125 <= pivot_out_3_124;
         start_in_3_125 <= start_out_3_124;
         swap_in_3_125 <= swap_out_3_124;
     end

     always @(posedge clk) begin
         data_in_3_125 <= data_out_2_125;
     end
  
     processor_AB AB_3_125 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_125),
       .start_in   (start_in_3_125),
       .swap_in   (swap_in_3_125),
       .op_in      (op_in_3_125),
       .pivot_in   (pivot_in_3_125),
       .start_out  (start_out_3_125),
       .swap_out   (swap_out_3_125),
       .data_out   (data_out_3_125),
       .op_out     (op_out_3_125),
       .pivot_out  (pivot_out_3_125),
       .r          (r_3_125)
     );

  // row 3, col 126

     reg start_in_3_126;
     wire start_out_3_126;

     reg swap_in_3_126;
     wire swap_out_3_126;

     reg [1:0] op_in_3_126;
     wire [1:0] op_out_3_126;

     wire r_3_126;

     reg data_in_3_126;
     wire data_out_3_126;

     reg pivot_in_3_126;
     wire pivot_out_3_126;

     always @(posedge clk) begin
         op_in_3_126 <= op_out_3_125;
         pivot_in_3_126 <= pivot_out_3_125;
         start_in_3_126 <= start_out_3_125;
         swap_in_3_126 <= swap_out_3_125;
     end

     always @(posedge clk) begin
         data_in_3_126 <= data_out_2_126;
     end
  
     processor_AB AB_3_126 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_126),
       .start_in   (start_in_3_126),
       .swap_in   (swap_in_3_126),
       .op_in      (op_in_3_126),
       .pivot_in   (pivot_in_3_126),
       .start_out  (start_out_3_126),
       .swap_out   (swap_out_3_126),
       .data_out   (data_out_3_126),
       .op_out     (op_out_3_126),
       .pivot_out  (pivot_out_3_126),
       .r          (r_3_126)
     );

  // row 3, col 127

     reg start_in_3_127;
     wire start_out_3_127;

     reg swap_in_3_127;
     wire swap_out_3_127;

     reg [1:0] op_in_3_127;
     wire [1:0] op_out_3_127;

     wire r_3_127;

     reg data_in_3_127;
     wire data_out_3_127;

     reg pivot_in_3_127;
     wire pivot_out_3_127;

     always @(posedge clk) begin
         op_in_3_127 <= op_out_3_126;
         pivot_in_3_127 <= pivot_out_3_126;
         start_in_3_127 <= start_out_3_126;
         swap_in_3_127 <= swap_out_3_126;
     end

     always @(posedge clk) begin
         data_in_3_127 <= data_out_2_127;
     end
  
     processor_AB AB_3_127 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_127),
       .start_in   (start_in_3_127),
       .swap_in   (swap_in_3_127),
       .op_in      (op_in_3_127),
       .pivot_in   (pivot_in_3_127),
       .start_out  (start_out_3_127),
       .swap_out   (swap_out_3_127),
       .data_out   (data_out_3_127),
       .op_out     (op_out_3_127),
       .pivot_out  (pivot_out_3_127),
       .r          (r_3_127)
     );

  // row 3, col 128

     reg start_in_3_128;
     wire start_out_3_128;

     reg swap_in_3_128;
     wire swap_out_3_128;

     reg [1:0] op_in_3_128;
     wire [1:0] op_out_3_128;

     wire r_3_128;

     reg data_in_3_128;
     wire data_out_3_128;

     reg pivot_in_3_128;
     wire pivot_out_3_128;

     always @(posedge clk) begin
         op_in_3_128 <= op_out_3_127;
         pivot_in_3_128 <= pivot_out_3_127;
         start_in_3_128 <= start_out_3_127;
         swap_in_3_128 <= swap_out_3_127;
     end

     always @(posedge clk) begin
         data_in_3_128 <= data_out_2_128;
     end
  
     processor_AB AB_3_128 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_128),
       .start_in   (start_in_3_128),
       .swap_in   (swap_in_3_128),
       .op_in      (op_in_3_128),
       .pivot_in   (pivot_in_3_128),
       .start_out  (start_out_3_128),
       .swap_out   (swap_out_3_128),
       .data_out   (data_out_3_128),
       .op_out     (op_out_3_128),
       .pivot_out  (pivot_out_3_128),
       .r          (r_3_128)
     );

  // row 3, col 129

     reg start_in_3_129;
     wire start_out_3_129;

     reg swap_in_3_129;
     wire swap_out_3_129;

     reg [1:0] op_in_3_129;
     wire [1:0] op_out_3_129;

     wire r_3_129;

     reg data_in_3_129;
     wire data_out_3_129;

     reg pivot_in_3_129;
     wire pivot_out_3_129;

     always @(posedge clk) begin
         op_in_3_129 <= op_out_3_128;
         pivot_in_3_129 <= pivot_out_3_128;
         start_in_3_129 <= start_out_3_128;
         swap_in_3_129 <= swap_out_3_128;
     end

     always @(posedge clk) begin
         data_in_3_129 <= data_out_2_129;
     end
  
     processor_AB AB_3_129 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_129),
       .start_in   (start_in_3_129),
       .swap_in   (swap_in_3_129),
       .op_in      (op_in_3_129),
       .pivot_in   (pivot_in_3_129),
       .start_out  (start_out_3_129),
       .swap_out   (swap_out_3_129),
       .data_out   (data_out_3_129),
       .op_out     (op_out_3_129),
       .pivot_out  (pivot_out_3_129),
       .r          (r_3_129)
     );

  // row 3, col 130

     reg start_in_3_130;
     wire start_out_3_130;

     reg swap_in_3_130;
     wire swap_out_3_130;

     reg [1:0] op_in_3_130;
     wire [1:0] op_out_3_130;

     wire r_3_130;

     reg data_in_3_130;
     wire data_out_3_130;

     reg pivot_in_3_130;
     wire pivot_out_3_130;

     always @(posedge clk) begin
         op_in_3_130 <= op_out_3_129;
         pivot_in_3_130 <= pivot_out_3_129;
         start_in_3_130 <= start_out_3_129;
         swap_in_3_130 <= swap_out_3_129;
     end

     always @(posedge clk) begin
         data_in_3_130 <= data_out_2_130;
     end
  
     processor_AB AB_3_130 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_130),
       .start_in   (start_in_3_130),
       .swap_in   (swap_in_3_130),
       .op_in      (op_in_3_130),
       .pivot_in   (pivot_in_3_130),
       .start_out  (start_out_3_130),
       .swap_out   (swap_out_3_130),
       .data_out   (data_out_3_130),
       .op_out     (op_out_3_130),
       .pivot_out  (pivot_out_3_130),
       .r          (r_3_130)
     );

  // row 3, col 131

     reg start_in_3_131;
     wire start_out_3_131;

     reg swap_in_3_131;
     wire swap_out_3_131;

     reg [1:0] op_in_3_131;
     wire [1:0] op_out_3_131;

     wire r_3_131;

     reg data_in_3_131;
     wire data_out_3_131;

     reg pivot_in_3_131;
     wire pivot_out_3_131;

     always @(posedge clk) begin
         op_in_3_131 <= op_out_3_130;
         pivot_in_3_131 <= pivot_out_3_130;
         start_in_3_131 <= start_out_3_130;
         swap_in_3_131 <= swap_out_3_130;
     end

     always @(posedge clk) begin
         data_in_3_131 <= data_out_2_131;
     end
  
     processor_AB AB_3_131 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_131),
       .start_in   (start_in_3_131),
       .swap_in   (swap_in_3_131),
       .op_in      (op_in_3_131),
       .pivot_in   (pivot_in_3_131),
       .start_out  (start_out_3_131),
       .swap_out   (swap_out_3_131),
       .data_out   (data_out_3_131),
       .op_out     (op_out_3_131),
       .pivot_out  (pivot_out_3_131),
       .r          (r_3_131)
     );

  // row 3, col 132

     reg start_in_3_132;
     wire start_out_3_132;

     reg swap_in_3_132;
     wire swap_out_3_132;

     reg [1:0] op_in_3_132;
     wire [1:0] op_out_3_132;

     wire r_3_132;

     reg data_in_3_132;
     wire data_out_3_132;

     reg pivot_in_3_132;
     wire pivot_out_3_132;

     always @(posedge clk) begin
         op_in_3_132 <= op_out_3_131;
         pivot_in_3_132 <= pivot_out_3_131;
         start_in_3_132 <= start_out_3_131;
         swap_in_3_132 <= swap_out_3_131;
     end

     always @(posedge clk) begin
         data_in_3_132 <= data_out_2_132;
     end
  
     processor_AB AB_3_132 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_132),
       .start_in   (start_in_3_132),
       .swap_in   (swap_in_3_132),
       .op_in      (op_in_3_132),
       .pivot_in   (pivot_in_3_132),
       .start_out  (start_out_3_132),
       .swap_out   (swap_out_3_132),
       .data_out   (data_out_3_132),
       .op_out     (op_out_3_132),
       .pivot_out  (pivot_out_3_132),
       .r          (r_3_132)
     );

  // row 3, col 133

     reg start_in_3_133;
     wire start_out_3_133;

     reg swap_in_3_133;
     wire swap_out_3_133;

     reg [1:0] op_in_3_133;
     wire [1:0] op_out_3_133;

     wire r_3_133;

     reg data_in_3_133;
     wire data_out_3_133;

     reg pivot_in_3_133;
     wire pivot_out_3_133;

     always @(posedge clk) begin
         op_in_3_133 <= op_out_3_132;
         pivot_in_3_133 <= pivot_out_3_132;
         start_in_3_133 <= start_out_3_132;
         swap_in_3_133 <= swap_out_3_132;
     end

     always @(posedge clk) begin
         data_in_3_133 <= data_out_2_133;
     end
  
     processor_AB AB_3_133 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_133),
       .start_in   (start_in_3_133),
       .swap_in   (swap_in_3_133),
       .op_in      (op_in_3_133),
       .pivot_in   (pivot_in_3_133),
       .start_out  (start_out_3_133),
       .swap_out   (swap_out_3_133),
       .data_out   (data_out_3_133),
       .op_out     (op_out_3_133),
       .pivot_out  (pivot_out_3_133),
       .r          (r_3_133)
     );

  // row 3, col 134

     reg start_in_3_134;
     wire start_out_3_134;

     reg swap_in_3_134;
     wire swap_out_3_134;

     reg [1:0] op_in_3_134;
     wire [1:0] op_out_3_134;

     wire r_3_134;

     reg data_in_3_134;
     wire data_out_3_134;

     reg pivot_in_3_134;
     wire pivot_out_3_134;

     always @(posedge clk) begin
         op_in_3_134 <= op_out_3_133;
         pivot_in_3_134 <= pivot_out_3_133;
         start_in_3_134 <= start_out_3_133;
         swap_in_3_134 <= swap_out_3_133;
     end

     always @(posedge clk) begin
         data_in_3_134 <= data_out_2_134;
     end
  
     processor_AB AB_3_134 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_134),
       .start_in   (start_in_3_134),
       .swap_in   (swap_in_3_134),
       .op_in      (op_in_3_134),
       .pivot_in   (pivot_in_3_134),
       .start_out  (start_out_3_134),
       .swap_out   (swap_out_3_134),
       .data_out   (data_out_3_134),
       .op_out     (op_out_3_134),
       .pivot_out  (pivot_out_3_134),
       .r          (r_3_134)
     );

  // row 3, col 135

     reg start_in_3_135;
     wire start_out_3_135;

     reg swap_in_3_135;
     wire swap_out_3_135;

     reg [1:0] op_in_3_135;
     wire [1:0] op_out_3_135;

     wire r_3_135;

     reg data_in_3_135;
     wire data_out_3_135;

     reg pivot_in_3_135;
     wire pivot_out_3_135;

     always @(posedge clk) begin
         op_in_3_135 <= op_out_3_134;
         pivot_in_3_135 <= pivot_out_3_134;
         start_in_3_135 <= start_out_3_134;
         swap_in_3_135 <= swap_out_3_134;
     end

     always @(posedge clk) begin
         data_in_3_135 <= data_out_2_135;
     end
  
     processor_AB AB_3_135 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_135),
       .start_in   (start_in_3_135),
       .swap_in   (swap_in_3_135),
       .op_in      (op_in_3_135),
       .pivot_in   (pivot_in_3_135),
       .start_out  (start_out_3_135),
       .swap_out   (swap_out_3_135),
       .data_out   (data_out_3_135),
       .op_out     (op_out_3_135),
       .pivot_out  (pivot_out_3_135),
       .r          (r_3_135)
     );

  // row 3, col 136

     reg start_in_3_136;
     wire start_out_3_136;

     reg swap_in_3_136;
     wire swap_out_3_136;

     reg [1:0] op_in_3_136;
     wire [1:0] op_out_3_136;

     wire r_3_136;

     reg data_in_3_136;
     wire data_out_3_136;

     reg pivot_in_3_136;
     wire pivot_out_3_136;

     always @(posedge clk) begin
         op_in_3_136 <= op_out_3_135;
         pivot_in_3_136 <= pivot_out_3_135;
         start_in_3_136 <= start_out_3_135;
         swap_in_3_136 <= swap_out_3_135;
     end

     always @(posedge clk) begin
         data_in_3_136 <= data_out_2_136;
     end
  
     processor_AB AB_3_136 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_136),
       .start_in   (start_in_3_136),
       .swap_in   (swap_in_3_136),
       .op_in      (op_in_3_136),
       .pivot_in   (pivot_in_3_136),
       .start_out  (start_out_3_136),
       .swap_out   (swap_out_3_136),
       .data_out   (data_out_3_136),
       .op_out     (op_out_3_136),
       .pivot_out  (pivot_out_3_136),
       .r          (r_3_136)
     );

  // row 3, col 137

     reg start_in_3_137;
     wire start_out_3_137;

     reg swap_in_3_137;
     wire swap_out_3_137;

     reg [1:0] op_in_3_137;
     wire [1:0] op_out_3_137;

     wire r_3_137;

     reg data_in_3_137;
     wire data_out_3_137;

     reg pivot_in_3_137;
     wire pivot_out_3_137;

     always @(posedge clk) begin
         op_in_3_137 <= op_out_3_136;
         pivot_in_3_137 <= pivot_out_3_136;
         start_in_3_137 <= start_out_3_136;
         swap_in_3_137 <= swap_out_3_136;
     end

     always @(posedge clk) begin
         data_in_3_137 <= data_out_2_137;
     end
  
     processor_AB AB_3_137 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_137),
       .start_in   (start_in_3_137),
       .swap_in   (swap_in_3_137),
       .op_in      (op_in_3_137),
       .pivot_in   (pivot_in_3_137),
       .start_out  (start_out_3_137),
       .swap_out   (swap_out_3_137),
       .data_out   (data_out_3_137),
       .op_out     (op_out_3_137),
       .pivot_out  (pivot_out_3_137),
       .r          (r_3_137)
     );

  // row 3, col 138

     reg start_in_3_138;
     wire start_out_3_138;

     reg swap_in_3_138;
     wire swap_out_3_138;

     reg [1:0] op_in_3_138;
     wire [1:0] op_out_3_138;

     wire r_3_138;

     reg data_in_3_138;
     wire data_out_3_138;

     reg pivot_in_3_138;
     wire pivot_out_3_138;

     always @(posedge clk) begin
         op_in_3_138 <= op_out_3_137;
         pivot_in_3_138 <= pivot_out_3_137;
         start_in_3_138 <= start_out_3_137;
         swap_in_3_138 <= swap_out_3_137;
     end

     always @(posedge clk) begin
         data_in_3_138 <= data_out_2_138;
     end
  
     processor_AB AB_3_138 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_138),
       .start_in   (start_in_3_138),
       .swap_in   (swap_in_3_138),
       .op_in      (op_in_3_138),
       .pivot_in   (pivot_in_3_138),
       .start_out  (start_out_3_138),
       .swap_out   (swap_out_3_138),
       .data_out   (data_out_3_138),
       .op_out     (op_out_3_138),
       .pivot_out  (pivot_out_3_138),
       .r          (r_3_138)
     );

  // row 3, col 139

     reg start_in_3_139;
     wire start_out_3_139;

     reg swap_in_3_139;
     wire swap_out_3_139;

     reg [1:0] op_in_3_139;
     wire [1:0] op_out_3_139;

     wire r_3_139;

     reg data_in_3_139;
     wire data_out_3_139;

     reg pivot_in_3_139;
     wire pivot_out_3_139;

     always @(posedge clk) begin
         op_in_3_139 <= op_out_3_138;
         pivot_in_3_139 <= pivot_out_3_138;
         start_in_3_139 <= start_out_3_138;
         swap_in_3_139 <= swap_out_3_138;
     end

     always @(posedge clk) begin
         data_in_3_139 <= data_out_2_139;
     end
  
     processor_AB AB_3_139 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_139),
       .start_in   (start_in_3_139),
       .swap_in   (swap_in_3_139),
       .op_in      (op_in_3_139),
       .pivot_in   (pivot_in_3_139),
       .start_out  (start_out_3_139),
       .swap_out   (swap_out_3_139),
       .data_out   (data_out_3_139),
       .op_out     (op_out_3_139),
       .pivot_out  (pivot_out_3_139),
       .r          (r_3_139)
     );

  // row 3, col 140

     reg start_in_3_140;
     wire start_out_3_140;

     reg swap_in_3_140;
     wire swap_out_3_140;

     reg [1:0] op_in_3_140;
     wire [1:0] op_out_3_140;

     wire r_3_140;

     reg data_in_3_140;
     wire data_out_3_140;

     reg pivot_in_3_140;
     wire pivot_out_3_140;

     always @(posedge clk) begin
         op_in_3_140 <= op_out_3_139;
         pivot_in_3_140 <= pivot_out_3_139;
         start_in_3_140 <= start_out_3_139;
         swap_in_3_140 <= swap_out_3_139;
     end

     always @(posedge clk) begin
         data_in_3_140 <= data_out_2_140;
     end
  
     processor_AB AB_3_140 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_140),
       .start_in   (start_in_3_140),
       .swap_in   (swap_in_3_140),
       .op_in      (op_in_3_140),
       .pivot_in   (pivot_in_3_140),
       .start_out  (start_out_3_140),
       .swap_out   (swap_out_3_140),
       .data_out   (data_out_3_140),
       .op_out     (op_out_3_140),
       .pivot_out  (pivot_out_3_140),
       .r          (r_3_140)
     );

  // row 3, col 141

     reg start_in_3_141;
     wire start_out_3_141;

     reg swap_in_3_141;
     wire swap_out_3_141;

     reg [1:0] op_in_3_141;
     wire [1:0] op_out_3_141;

     wire r_3_141;

     reg data_in_3_141;
     wire data_out_3_141;

     reg pivot_in_3_141;
     wire pivot_out_3_141;

     always @(posedge clk) begin
         op_in_3_141 <= op_out_3_140;
         pivot_in_3_141 <= pivot_out_3_140;
         start_in_3_141 <= start_out_3_140;
         swap_in_3_141 <= swap_out_3_140;
     end

     always @(posedge clk) begin
         data_in_3_141 <= data_out_2_141;
     end
  
     processor_AB AB_3_141 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_141),
       .start_in   (start_in_3_141),
       .swap_in   (swap_in_3_141),
       .op_in      (op_in_3_141),
       .pivot_in   (pivot_in_3_141),
       .start_out  (start_out_3_141),
       .swap_out   (swap_out_3_141),
       .data_out   (data_out_3_141),
       .op_out     (op_out_3_141),
       .pivot_out  (pivot_out_3_141),
       .r          (r_3_141)
     );

  // row 3, col 142

     reg start_in_3_142;
     wire start_out_3_142;

     reg swap_in_3_142;
     wire swap_out_3_142;

     reg [1:0] op_in_3_142;
     wire [1:0] op_out_3_142;

     wire r_3_142;

     reg data_in_3_142;
     wire data_out_3_142;

     reg pivot_in_3_142;
     wire pivot_out_3_142;

     always @(posedge clk) begin
         op_in_3_142 <= op_out_3_141;
         pivot_in_3_142 <= pivot_out_3_141;
         start_in_3_142 <= start_out_3_141;
         swap_in_3_142 <= swap_out_3_141;
     end

     always @(posedge clk) begin
         data_in_3_142 <= data_out_2_142;
     end
  
     processor_AB AB_3_142 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_142),
       .start_in   (start_in_3_142),
       .swap_in   (swap_in_3_142),
       .op_in      (op_in_3_142),
       .pivot_in   (pivot_in_3_142),
       .start_out  (start_out_3_142),
       .swap_out   (swap_out_3_142),
       .data_out   (data_out_3_142),
       .op_out     (op_out_3_142),
       .pivot_out  (pivot_out_3_142),
       .r          (r_3_142)
     );

  // row 3, col 143

     reg start_in_3_143;
     wire start_out_3_143;

     reg swap_in_3_143;
     wire swap_out_3_143;

     reg [1:0] op_in_3_143;
     wire [1:0] op_out_3_143;

     wire r_3_143;

     reg data_in_3_143;
     wire data_out_3_143;

     reg pivot_in_3_143;
     wire pivot_out_3_143;

     always @(posedge clk) begin
         op_in_3_143 <= op_out_3_142;
         pivot_in_3_143 <= pivot_out_3_142;
         start_in_3_143 <= start_out_3_142;
         swap_in_3_143 <= swap_out_3_142;
     end

     always @(posedge clk) begin
         data_in_3_143 <= data_out_2_143;
     end
  
     processor_AB AB_3_143 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_143),
       .start_in   (start_in_3_143),
       .swap_in   (swap_in_3_143),
       .op_in      (op_in_3_143),
       .pivot_in   (pivot_in_3_143),
       .start_out  (start_out_3_143),
       .swap_out   (swap_out_3_143),
       .data_out   (data_out_3_143),
       .op_out     (op_out_3_143),
       .pivot_out  (pivot_out_3_143),
       .r          (r_3_143)
     );

  // row 3, col 144

     reg start_in_3_144;
     wire start_out_3_144;

     reg swap_in_3_144;
     wire swap_out_3_144;

     reg [1:0] op_in_3_144;
     wire [1:0] op_out_3_144;

     wire r_3_144;

     reg data_in_3_144;
     wire data_out_3_144;

     reg pivot_in_3_144;
     wire pivot_out_3_144;

     always @(posedge clk) begin
         op_in_3_144 <= op_out_3_143;
         pivot_in_3_144 <= pivot_out_3_143;
         start_in_3_144 <= start_out_3_143;
         swap_in_3_144 <= swap_out_3_143;
     end

     always @(posedge clk) begin
         data_in_3_144 <= data_out_2_144;
     end
  
     processor_AB AB_3_144 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_144),
       .start_in   (start_in_3_144),
       .swap_in   (swap_in_3_144),
       .op_in      (op_in_3_144),
       .pivot_in   (pivot_in_3_144),
       .start_out  (start_out_3_144),
       .swap_out   (swap_out_3_144),
       .data_out   (data_out_3_144),
       .op_out     (op_out_3_144),
       .pivot_out  (pivot_out_3_144),
       .r          (r_3_144)
     );

  // row 3, col 145

     reg start_in_3_145;
     wire start_out_3_145;

     reg swap_in_3_145;
     wire swap_out_3_145;

     reg [1:0] op_in_3_145;
     wire [1:0] op_out_3_145;

     wire r_3_145;

     reg data_in_3_145;
     wire data_out_3_145;

     reg pivot_in_3_145;
     wire pivot_out_3_145;

     always @(posedge clk) begin
         op_in_3_145 <= op_out_3_144;
         pivot_in_3_145 <= pivot_out_3_144;
         start_in_3_145 <= start_out_3_144;
         swap_in_3_145 <= swap_out_3_144;
     end

     always @(posedge clk) begin
         data_in_3_145 <= data_out_2_145;
     end
  
     processor_AB AB_3_145 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_145),
       .start_in   (start_in_3_145),
       .swap_in   (swap_in_3_145),
       .op_in      (op_in_3_145),
       .pivot_in   (pivot_in_3_145),
       .start_out  (start_out_3_145),
       .swap_out   (swap_out_3_145),
       .data_out   (data_out_3_145),
       .op_out     (op_out_3_145),
       .pivot_out  (pivot_out_3_145),
       .r          (r_3_145)
     );

  // row 3, col 146

     reg start_in_3_146;
     wire start_out_3_146;

     reg swap_in_3_146;
     wire swap_out_3_146;

     reg [1:0] op_in_3_146;
     wire [1:0] op_out_3_146;

     wire r_3_146;

     reg data_in_3_146;
     wire data_out_3_146;

     reg pivot_in_3_146;
     wire pivot_out_3_146;

     always @(posedge clk) begin
         op_in_3_146 <= op_out_3_145;
         pivot_in_3_146 <= pivot_out_3_145;
         start_in_3_146 <= start_out_3_145;
         swap_in_3_146 <= swap_out_3_145;
     end

     always @(posedge clk) begin
         data_in_3_146 <= data_out_2_146;
     end
  
     processor_AB AB_3_146 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_146),
       .start_in   (start_in_3_146),
       .swap_in   (swap_in_3_146),
       .op_in      (op_in_3_146),
       .pivot_in   (pivot_in_3_146),
       .start_out  (start_out_3_146),
       .swap_out   (swap_out_3_146),
       .data_out   (data_out_3_146),
       .op_out     (op_out_3_146),
       .pivot_out  (pivot_out_3_146),
       .r          (r_3_146)
     );

  // row 3, col 147

     reg start_in_3_147;
     wire start_out_3_147;

     reg swap_in_3_147;
     wire swap_out_3_147;

     reg [1:0] op_in_3_147;
     wire [1:0] op_out_3_147;

     wire r_3_147;

     reg data_in_3_147;
     wire data_out_3_147;

     reg pivot_in_3_147;
     wire pivot_out_3_147;

     always @(posedge clk) begin
         op_in_3_147 <= op_out_3_146;
         pivot_in_3_147 <= pivot_out_3_146;
         start_in_3_147 <= start_out_3_146;
         swap_in_3_147 <= swap_out_3_146;
     end

     always @(posedge clk) begin
         data_in_3_147 <= data_out_2_147;
     end
  
     processor_AB AB_3_147 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_147),
       .start_in   (start_in_3_147),
       .swap_in   (swap_in_3_147),
       .op_in      (op_in_3_147),
       .pivot_in   (pivot_in_3_147),
       .start_out  (start_out_3_147),
       .swap_out   (swap_out_3_147),
       .data_out   (data_out_3_147),
       .op_out     (op_out_3_147),
       .pivot_out  (pivot_out_3_147),
       .r          (r_3_147)
     );

  // row 3, col 148

     reg start_in_3_148;
     wire start_out_3_148;

     reg swap_in_3_148;
     wire swap_out_3_148;

     reg [1:0] op_in_3_148;
     wire [1:0] op_out_3_148;

     wire r_3_148;

     reg data_in_3_148;
     wire data_out_3_148;

     reg pivot_in_3_148;
     wire pivot_out_3_148;

     always @(posedge clk) begin
         op_in_3_148 <= op_out_3_147;
         pivot_in_3_148 <= pivot_out_3_147;
         start_in_3_148 <= start_out_3_147;
         swap_in_3_148 <= swap_out_3_147;
     end

     always @(posedge clk) begin
         data_in_3_148 <= data_out_2_148;
     end
  
     processor_AB AB_3_148 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_148),
       .start_in   (start_in_3_148),
       .swap_in   (swap_in_3_148),
       .op_in      (op_in_3_148),
       .pivot_in   (pivot_in_3_148),
       .start_out  (start_out_3_148),
       .swap_out   (swap_out_3_148),
       .data_out   (data_out_3_148),
       .op_out     (op_out_3_148),
       .pivot_out  (pivot_out_3_148),
       .r          (r_3_148)
     );

  // row 3, col 149

     reg start_in_3_149;
     wire start_out_3_149;

     reg swap_in_3_149;
     wire swap_out_3_149;

     reg [1:0] op_in_3_149;
     wire [1:0] op_out_3_149;

     wire r_3_149;

     reg data_in_3_149;
     wire data_out_3_149;

     reg pivot_in_3_149;
     wire pivot_out_3_149;

     always @(posedge clk) begin
         op_in_3_149 <= op_out_3_148;
         pivot_in_3_149 <= pivot_out_3_148;
         start_in_3_149 <= start_out_3_148;
         swap_in_3_149 <= swap_out_3_148;
     end

     always @(posedge clk) begin
         data_in_3_149 <= data_out_2_149;
     end
  
     processor_AB AB_3_149 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_149),
       .start_in   (start_in_3_149),
       .swap_in   (swap_in_3_149),
       .op_in      (op_in_3_149),
       .pivot_in   (pivot_in_3_149),
       .start_out  (start_out_3_149),
       .swap_out   (swap_out_3_149),
       .data_out   (data_out_3_149),
       .op_out     (op_out_3_149),
       .pivot_out  (pivot_out_3_149),
       .r          (r_3_149)
     );

  // row 3, col 150

     reg start_in_3_150;
     wire start_out_3_150;

     reg swap_in_3_150;
     wire swap_out_3_150;

     reg [1:0] op_in_3_150;
     wire [1:0] op_out_3_150;

     wire r_3_150;

     reg data_in_3_150;
     wire data_out_3_150;

     reg pivot_in_3_150;
     wire pivot_out_3_150;

     always @(posedge clk) begin
         op_in_3_150 <= op_out_3_149;
         pivot_in_3_150 <= pivot_out_3_149;
         start_in_3_150 <= start_out_3_149;
         swap_in_3_150 <= swap_out_3_149;
     end

     always @(posedge clk) begin
         data_in_3_150 <= data_out_2_150;
     end
  
     processor_AB AB_3_150 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_150),
       .start_in   (start_in_3_150),
       .swap_in   (swap_in_3_150),
       .op_in      (op_in_3_150),
       .pivot_in   (pivot_in_3_150),
       .start_out  (start_out_3_150),
       .swap_out   (swap_out_3_150),
       .data_out   (data_out_3_150),
       .op_out     (op_out_3_150),
       .pivot_out  (pivot_out_3_150),
       .r          (r_3_150)
     );

  // row 3, col 151

     reg start_in_3_151;
     wire start_out_3_151;

     reg swap_in_3_151;
     wire swap_out_3_151;

     reg [1:0] op_in_3_151;
     wire [1:0] op_out_3_151;

     wire r_3_151;

     reg data_in_3_151;
     wire data_out_3_151;

     reg pivot_in_3_151;
     wire pivot_out_3_151;

     always @(posedge clk) begin
         op_in_3_151 <= op_out_3_150;
         pivot_in_3_151 <= pivot_out_3_150;
         start_in_3_151 <= start_out_3_150;
         swap_in_3_151 <= swap_out_3_150;
     end

     always @(posedge clk) begin
         data_in_3_151 <= data_out_2_151;
     end
  
     processor_AB AB_3_151 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_151),
       .start_in   (start_in_3_151),
       .swap_in   (swap_in_3_151),
       .op_in      (op_in_3_151),
       .pivot_in   (pivot_in_3_151),
       .start_out  (start_out_3_151),
       .swap_out   (swap_out_3_151),
       .data_out   (data_out_3_151),
       .op_out     (op_out_3_151),
       .pivot_out  (pivot_out_3_151),
       .r          (r_3_151)
     );

  // row 3, col 152

     reg start_in_3_152;
     wire start_out_3_152;

     reg swap_in_3_152;
     wire swap_out_3_152;

     reg [1:0] op_in_3_152;
     wire [1:0] op_out_3_152;

     wire r_3_152;

     reg data_in_3_152;
     wire data_out_3_152;

     reg pivot_in_3_152;
     wire pivot_out_3_152;

     always @(posedge clk) begin
         op_in_3_152 <= op_out_3_151;
         pivot_in_3_152 <= pivot_out_3_151;
         start_in_3_152 <= start_out_3_151;
         swap_in_3_152 <= swap_out_3_151;
     end

     always @(posedge clk) begin
         data_in_3_152 <= data_out_2_152;
     end
  
     processor_AB AB_3_152 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_152),
       .start_in   (start_in_3_152),
       .swap_in   (swap_in_3_152),
       .op_in      (op_in_3_152),
       .pivot_in   (pivot_in_3_152),
       .start_out  (start_out_3_152),
       .swap_out   (swap_out_3_152),
       .data_out   (data_out_3_152),
       .op_out     (op_out_3_152),
       .pivot_out  (pivot_out_3_152),
       .r          (r_3_152)
     );

  // row 3, col 153

     reg start_in_3_153;
     wire start_out_3_153;

     reg swap_in_3_153;
     wire swap_out_3_153;

     reg [1:0] op_in_3_153;
     wire [1:0] op_out_3_153;

     wire r_3_153;

     reg data_in_3_153;
     wire data_out_3_153;

     reg pivot_in_3_153;
     wire pivot_out_3_153;

     always @(posedge clk) begin
         op_in_3_153 <= op_out_3_152;
         pivot_in_3_153 <= pivot_out_3_152;
         start_in_3_153 <= start_out_3_152;
         swap_in_3_153 <= swap_out_3_152;
     end

     always @(posedge clk) begin
         data_in_3_153 <= data_out_2_153;
     end
  
     processor_AB AB_3_153 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_153),
       .start_in   (start_in_3_153),
       .swap_in   (swap_in_3_153),
       .op_in      (op_in_3_153),
       .pivot_in   (pivot_in_3_153),
       .start_out  (start_out_3_153),
       .swap_out   (swap_out_3_153),
       .data_out   (data_out_3_153),
       .op_out     (op_out_3_153),
       .pivot_out  (pivot_out_3_153),
       .r          (r_3_153)
     );

  // row 3, col 154

     reg start_in_3_154;
     wire start_out_3_154;

     reg swap_in_3_154;
     wire swap_out_3_154;

     reg [1:0] op_in_3_154;
     wire [1:0] op_out_3_154;

     wire r_3_154;

     reg data_in_3_154;
     wire data_out_3_154;

     reg pivot_in_3_154;
     wire pivot_out_3_154;

     always @(posedge clk) begin
         op_in_3_154 <= op_out_3_153;
         pivot_in_3_154 <= pivot_out_3_153;
         start_in_3_154 <= start_out_3_153;
         swap_in_3_154 <= swap_out_3_153;
     end

     always @(posedge clk) begin
         data_in_3_154 <= data_out_2_154;
     end
  
     processor_AB AB_3_154 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_154),
       .start_in   (start_in_3_154),
       .swap_in   (swap_in_3_154),
       .op_in      (op_in_3_154),
       .pivot_in   (pivot_in_3_154),
       .start_out  (start_out_3_154),
       .swap_out   (swap_out_3_154),
       .data_out   (data_out_3_154),
       .op_out     (op_out_3_154),
       .pivot_out  (pivot_out_3_154),
       .r          (r_3_154)
     );

  // row 3, col 155

     reg start_in_3_155;
     wire start_out_3_155;

     reg swap_in_3_155;
     wire swap_out_3_155;

     reg [1:0] op_in_3_155;
     wire [1:0] op_out_3_155;

     wire r_3_155;

     reg data_in_3_155;
     wire data_out_3_155;

     reg pivot_in_3_155;
     wire pivot_out_3_155;

     always @(posedge clk) begin
         op_in_3_155 <= op_out_3_154;
         pivot_in_3_155 <= pivot_out_3_154;
         start_in_3_155 <= start_out_3_154;
         swap_in_3_155 <= swap_out_3_154;
     end

     always @(posedge clk) begin
         data_in_3_155 <= data_out_2_155;
     end
  
     processor_AB AB_3_155 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_155),
       .start_in   (start_in_3_155),
       .swap_in   (swap_in_3_155),
       .op_in      (op_in_3_155),
       .pivot_in   (pivot_in_3_155),
       .start_out  (start_out_3_155),
       .swap_out   (swap_out_3_155),
       .data_out   (data_out_3_155),
       .op_out     (op_out_3_155),
       .pivot_out  (pivot_out_3_155),
       .r          (r_3_155)
     );

  // row 3, col 156

     reg start_in_3_156;
     wire start_out_3_156;

     reg swap_in_3_156;
     wire swap_out_3_156;

     reg [1:0] op_in_3_156;
     wire [1:0] op_out_3_156;

     wire r_3_156;

     reg data_in_3_156;
     wire data_out_3_156;

     reg pivot_in_3_156;
     wire pivot_out_3_156;

     always @(posedge clk) begin
         op_in_3_156 <= op_out_3_155;
         pivot_in_3_156 <= pivot_out_3_155;
         start_in_3_156 <= start_out_3_155;
         swap_in_3_156 <= swap_out_3_155;
     end

     always @(posedge clk) begin
         data_in_3_156 <= data_out_2_156;
     end
  
     processor_AB AB_3_156 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_156),
       .start_in   (start_in_3_156),
       .swap_in   (swap_in_3_156),
       .op_in      (op_in_3_156),
       .pivot_in   (pivot_in_3_156),
       .start_out  (start_out_3_156),
       .swap_out   (swap_out_3_156),
       .data_out   (data_out_3_156),
       .op_out     (op_out_3_156),
       .pivot_out  (pivot_out_3_156),
       .r          (r_3_156)
     );

  // row 3, col 157

     reg start_in_3_157;
     wire start_out_3_157;

     reg swap_in_3_157;
     wire swap_out_3_157;

     reg [1:0] op_in_3_157;
     wire [1:0] op_out_3_157;

     wire r_3_157;

     reg data_in_3_157;
     wire data_out_3_157;

     reg pivot_in_3_157;
     wire pivot_out_3_157;

     always @(posedge clk) begin
         op_in_3_157 <= op_out_3_156;
         pivot_in_3_157 <= pivot_out_3_156;
         start_in_3_157 <= start_out_3_156;
         swap_in_3_157 <= swap_out_3_156;
     end

     always @(posedge clk) begin
         data_in_3_157 <= data_out_2_157;
     end
  
     processor_AB AB_3_157 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_157),
       .start_in   (start_in_3_157),
       .swap_in   (swap_in_3_157),
       .op_in      (op_in_3_157),
       .pivot_in   (pivot_in_3_157),
       .start_out  (start_out_3_157),
       .swap_out   (swap_out_3_157),
       .data_out   (data_out_3_157),
       .op_out     (op_out_3_157),
       .pivot_out  (pivot_out_3_157),
       .r          (r_3_157)
     );

  // row 3, col 158

     reg start_in_3_158;
     wire start_out_3_158;

     reg swap_in_3_158;
     wire swap_out_3_158;

     reg [1:0] op_in_3_158;
     wire [1:0] op_out_3_158;

     wire r_3_158;

     reg data_in_3_158;
     wire data_out_3_158;

     reg pivot_in_3_158;
     wire pivot_out_3_158;

     always @(posedge clk) begin
         op_in_3_158 <= op_out_3_157;
         pivot_in_3_158 <= pivot_out_3_157;
         start_in_3_158 <= start_out_3_157;
         swap_in_3_158 <= swap_out_3_157;
     end

     always @(posedge clk) begin
         data_in_3_158 <= data_out_2_158;
     end
  
     processor_AB AB_3_158 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_158),
       .start_in   (start_in_3_158),
       .swap_in   (swap_in_3_158),
       .op_in      (op_in_3_158),
       .pivot_in   (pivot_in_3_158),
       .start_out  (start_out_3_158),
       .swap_out   (swap_out_3_158),
       .data_out   (data_out_3_158),
       .op_out     (op_out_3_158),
       .pivot_out  (pivot_out_3_158),
       .r          (r_3_158)
     );

  // row 3, col 159

     reg start_in_3_159;
     wire start_out_3_159;

     reg swap_in_3_159;
     wire swap_out_3_159;

     reg [1:0] op_in_3_159;
     wire [1:0] op_out_3_159;

     wire r_3_159;

     reg data_in_3_159;
     wire data_out_3_159;

     reg pivot_in_3_159;
     wire pivot_out_3_159;

     always @(posedge clk) begin
         op_in_3_159 <= op_out_3_158;
         pivot_in_3_159 <= pivot_out_3_158;
         start_in_3_159 <= start_out_3_158;
         swap_in_3_159 <= swap_out_3_158;
     end

     always @(posedge clk) begin
         data_in_3_159 <= data_out_2_159;
     end
  
     processor_AB AB_3_159 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_159),
       .start_in   (start_in_3_159),
       .swap_in   (swap_in_3_159),
       .op_in      (op_in_3_159),
       .pivot_in   (pivot_in_3_159),
       .start_out  (start_out_3_159),
       .swap_out   (swap_out_3_159),
       .data_out   (data_out_3_159),
       .op_out     (op_out_3_159),
       .pivot_out  (pivot_out_3_159),
       .r          (r_3_159)
     );

  // row 3, col 160

     reg start_in_3_160;
     wire start_out_3_160;

     reg swap_in_3_160;
     wire swap_out_3_160;

     reg [1:0] op_in_3_160;
     wire [1:0] op_out_3_160;

     wire r_3_160;

     reg data_in_3_160;
     wire data_out_3_160;

     reg pivot_in_3_160;
     wire pivot_out_3_160;

     always @(posedge clk) begin
         op_in_3_160 <= op_out_3_159;
         pivot_in_3_160 <= pivot_out_3_159;
         start_in_3_160 <= start_out_3_159;
         swap_in_3_160 <= swap_out_3_159;
     end

     always @(posedge clk) begin
         data_in_3_160 <= data_out_2_160;
     end
  
     processor_AB AB_3_160 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_160),
       .start_in   (start_in_3_160),
       .swap_in   (swap_in_3_160),
       .op_in      (op_in_3_160),
       .pivot_in   (pivot_in_3_160),
       .start_out  (start_out_3_160),
       .swap_out   (swap_out_3_160),
       .data_out   (data_out_3_160),
       .op_out     (op_out_3_160),
       .pivot_out  (pivot_out_3_160),
       .r          (r_3_160)
     );

  // row 3, col 161

     reg start_in_3_161;
     wire start_out_3_161;

     reg swap_in_3_161;
     wire swap_out_3_161;

     reg [1:0] op_in_3_161;
     wire [1:0] op_out_3_161;

     wire r_3_161;

     reg data_in_3_161;
     wire data_out_3_161;

     reg pivot_in_3_161;
     wire pivot_out_3_161;

     always @(posedge clk) begin
         op_in_3_161 <= op_out_3_160;
         pivot_in_3_161 <= pivot_out_3_160;
         start_in_3_161 <= start_out_3_160;
         swap_in_3_161 <= swap_out_3_160;
     end

     always @(posedge clk) begin
         data_in_3_161 <= data_out_2_161;
     end
  
     processor_AB AB_3_161 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_161),
       .start_in   (start_in_3_161),
       .swap_in   (swap_in_3_161),
       .op_in      (op_in_3_161),
       .pivot_in   (pivot_in_3_161),
       .start_out  (start_out_3_161),
       .swap_out   (swap_out_3_161),
       .data_out   (data_out_3_161),
       .op_out     (op_out_3_161),
       .pivot_out  (pivot_out_3_161),
       .r          (r_3_161)
     );

  // row 3, col 162

     reg start_in_3_162;
     wire start_out_3_162;

     reg swap_in_3_162;
     wire swap_out_3_162;

     reg [1:0] op_in_3_162;
     wire [1:0] op_out_3_162;

     wire r_3_162;

     reg data_in_3_162;
     wire data_out_3_162;

     reg pivot_in_3_162;
     wire pivot_out_3_162;

     always @(posedge clk) begin
         op_in_3_162 <= op_out_3_161;
         pivot_in_3_162 <= pivot_out_3_161;
         start_in_3_162 <= start_out_3_161;
         swap_in_3_162 <= swap_out_3_161;
     end

     always @(posedge clk) begin
         data_in_3_162 <= data_out_2_162;
     end
  
     processor_AB AB_3_162 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_162),
       .start_in   (start_in_3_162),
       .swap_in   (swap_in_3_162),
       .op_in      (op_in_3_162),
       .pivot_in   (pivot_in_3_162),
       .start_out  (start_out_3_162),
       .swap_out   (swap_out_3_162),
       .data_out   (data_out_3_162),
       .op_out     (op_out_3_162),
       .pivot_out  (pivot_out_3_162),
       .r          (r_3_162)
     );

  // row 3, col 163

     reg start_in_3_163;
     wire start_out_3_163;

     reg swap_in_3_163;
     wire swap_out_3_163;

     reg [1:0] op_in_3_163;
     wire [1:0] op_out_3_163;

     wire r_3_163;

     reg data_in_3_163;
     wire data_out_3_163;

     reg pivot_in_3_163;
     wire pivot_out_3_163;

     always @(posedge clk) begin
         op_in_3_163 <= op_out_3_162;
         pivot_in_3_163 <= pivot_out_3_162;
         start_in_3_163 <= start_out_3_162;
         swap_in_3_163 <= swap_out_3_162;
     end

     always @(posedge clk) begin
         data_in_3_163 <= data_out_2_163;
     end
  
     processor_AB AB_3_163 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_163),
       .start_in   (start_in_3_163),
       .swap_in   (swap_in_3_163),
       .op_in      (op_in_3_163),
       .pivot_in   (pivot_in_3_163),
       .start_out  (start_out_3_163),
       .swap_out   (swap_out_3_163),
       .data_out   (data_out_3_163),
       .op_out     (op_out_3_163),
       .pivot_out  (pivot_out_3_163),
       .r          (r_3_163)
     );

  // row 3, col 164

     reg start_in_3_164;
     wire start_out_3_164;

     reg swap_in_3_164;
     wire swap_out_3_164;

     reg [1:0] op_in_3_164;
     wire [1:0] op_out_3_164;

     wire r_3_164;

     reg data_in_3_164;
     wire data_out_3_164;

     reg pivot_in_3_164;
     wire pivot_out_3_164;

     always @(posedge clk) begin
         op_in_3_164 <= op_out_3_163;
         pivot_in_3_164 <= pivot_out_3_163;
         start_in_3_164 <= start_out_3_163;
         swap_in_3_164 <= swap_out_3_163;
     end

     always @(posedge clk) begin
         data_in_3_164 <= data_out_2_164;
     end
  
     processor_AB AB_3_164 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_164),
       .start_in   (start_in_3_164),
       .swap_in   (swap_in_3_164),
       .op_in      (op_in_3_164),
       .pivot_in   (pivot_in_3_164),
       .start_out  (start_out_3_164),
       .swap_out   (swap_out_3_164),
       .data_out   (data_out_3_164),
       .op_out     (op_out_3_164),
       .pivot_out  (pivot_out_3_164),
       .r          (r_3_164)
     );

  // row 3, col 165

     reg start_in_3_165;
     wire start_out_3_165;

     reg swap_in_3_165;
     wire swap_out_3_165;

     reg [1:0] op_in_3_165;
     wire [1:0] op_out_3_165;

     wire r_3_165;

     reg data_in_3_165;
     wire data_out_3_165;

     reg pivot_in_3_165;
     wire pivot_out_3_165;

     always @(posedge clk) begin
         op_in_3_165 <= op_out_3_164;
         pivot_in_3_165 <= pivot_out_3_164;
         start_in_3_165 <= start_out_3_164;
         swap_in_3_165 <= swap_out_3_164;
     end

     always @(posedge clk) begin
         data_in_3_165 <= data_out_2_165;
     end
  
     processor_AB AB_3_165 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_3_165),
       .start_in   (start_in_3_165),
       .swap_in   (swap_in_3_165),
       .op_in      (op_in_3_165),
       .pivot_in   (pivot_in_3_165),
       .start_out  (start_out_3_165),
       .swap_out   (swap_out_3_165),
       .data_out   (data_out_3_165),
       .op_out     (op_out_3_165),
       .pivot_out  (pivot_out_3_165),
       .r          (r_3_165)
     );

  /////////////////////////////////////
  // row 4
  // row 4, col 0

     wire start_in_4_0;
     wire start_out_4_0;

     wire swap_in_4_0;
     wire swap_out_4_0;

     wire [1:0] op_in_4_0;
     wire [1:0] op_out_4_0;

     wire r_4_0;

     reg data_in_4_0;
     wire data_out_4_0;

     wire pivot_in_4_0;
     wire pivout_out_4_0;

     assign op_in_4_0 = 2'b00;
     assign pivot_in_4_0 = 0;

     assign start_in_4_0 = start_row[4]; 
     assign swap_in_4_0 = mode ? swap : swap_row[4]; 

     always @(posedge clk) begin
         data_in_4_0 <= data_out_3_0;
     end

     processor_AB AB_4_0 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_0),
       .start_in   (start_in_4_0),
       .swap_in   (swap_in_4_0),
       .op_in      (op_in_4_0),
       .pivot_in   (pivot_in_4_0),
       .start_out  (start_out_4_0),
       .swap_out   (swap_out_4_0),
       .data_out   (data_out_4_0),
       .op_out     (op_out_4_0),
       .pivot_out  (pivot_out_4_0),
       .r          (r_4_0)
     );

  // row 4, col 1

     reg start_in_4_1;
     wire start_out_4_1;

     reg swap_in_4_1;
     wire swap_out_4_1;

     reg [1:0] op_in_4_1;
     wire [1:0] op_out_4_1;

     wire r_4_1;

     reg data_in_4_1;
     wire data_out_4_1;

     reg pivot_in_4_1;
     wire pivot_out_4_1;

     always @(posedge clk) begin
         op_in_4_1 <= op_out_4_0;
         pivot_in_4_1 <= pivot_out_4_0;
         start_in_4_1 <= start_out_4_0;
         swap_in_4_1 <= swap_out_4_0;
     end

     always @(posedge clk) begin
         data_in_4_1 <= data_out_3_1;
     end
  
     processor_AB AB_4_1 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_1),
       .start_in   (start_in_4_1),
       .swap_in   (swap_in_4_1),
       .op_in      (op_in_4_1),
       .pivot_in   (pivot_in_4_1),
       .start_out  (start_out_4_1),
       .swap_out   (swap_out_4_1),
       .data_out   (data_out_4_1),
       .op_out     (op_out_4_1),
       .pivot_out  (pivot_out_4_1),
       .r          (r_4_1)
     );

  // row 4, col 2

     reg start_in_4_2;
     wire start_out_4_2;

     reg swap_in_4_2;
     wire swap_out_4_2;

     reg [1:0] op_in_4_2;
     wire [1:0] op_out_4_2;

     wire r_4_2;

     reg data_in_4_2;
     wire data_out_4_2;

     reg pivot_in_4_2;
     wire pivot_out_4_2;

     always @(posedge clk) begin
         op_in_4_2 <= op_out_4_1;
         pivot_in_4_2 <= pivot_out_4_1;
         start_in_4_2 <= start_out_4_1;
         swap_in_4_2 <= swap_out_4_1;
     end

     always @(posedge clk) begin
         data_in_4_2 <= data_out_3_2;
     end
  
     processor_AB AB_4_2 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_2),
       .start_in   (start_in_4_2),
       .swap_in   (swap_in_4_2),
       .op_in      (op_in_4_2),
       .pivot_in   (pivot_in_4_2),
       .start_out  (start_out_4_2),
       .swap_out   (swap_out_4_2),
       .data_out   (data_out_4_2),
       .op_out     (op_out_4_2),
       .pivot_out  (pivot_out_4_2),
       .r          (r_4_2)
     );

  // row 4, col 3

     reg start_in_4_3;
     wire start_out_4_3;

     reg swap_in_4_3;
     wire swap_out_4_3;

     reg [1:0] op_in_4_3;
     wire [1:0] op_out_4_3;

     wire r_4_3;

     reg data_in_4_3;
     wire data_out_4_3;

     reg pivot_in_4_3;
     wire pivot_out_4_3;

     always @(posedge clk) begin
         op_in_4_3 <= op_out_4_2;
         pivot_in_4_3 <= pivot_out_4_2;
         start_in_4_3 <= start_out_4_2;
         swap_in_4_3 <= swap_out_4_2;
     end

     always @(posedge clk) begin
         data_in_4_3 <= data_out_3_3;
     end
  
     processor_AB AB_4_3 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_3),
       .start_in   (start_in_4_3),
       .swap_in   (swap_in_4_3),
       .op_in      (op_in_4_3),
       .pivot_in   (pivot_in_4_3),
       .start_out  (start_out_4_3),
       .swap_out   (swap_out_4_3),
       .data_out   (data_out_4_3),
       .op_out     (op_out_4_3),
       .pivot_out  (pivot_out_4_3),
       .r          (r_4_3)
     );

  // row 4, col 4

     reg start_in_4_4;
     wire start_out_4_4;

     reg swap_in_4_4;
     wire swap_out_4_4;

     reg [1:0] op_in_4_4;
     wire [1:0] op_out_4_4;

     wire r_4_4;

     reg data_in_4_4;
     wire data_out_4_4;

     reg pivot_in_4_4;
     wire pivot_out_4_4;

     always @(posedge clk) begin
         op_in_4_4 <= op_out_4_3;
         pivot_in_4_4 <= pivot_out_4_3;
         start_in_4_4 <= start_out_4_3;
         swap_in_4_4 <= swap_out_4_3;
     end

     always @(posedge clk) begin
         data_in_4_4 <= data_out_3_4;
     end
  
     processor_AB AB_4_4 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_4),
       .start_in   (start_in_4_4),
       .swap_in   (swap_in_4_4),
       .op_in      (op_in_4_4),
       .pivot_in   (pivot_in_4_4),
       .start_out  (start_out_4_4),
       .swap_out   (swap_out_4_4),
       .data_out   (data_out_4_4),
       .op_out     (op_out_4_4),
       .pivot_out  (pivot_out_4_4),
       .r          (r_4_4)
     );

  // row 4, col 5

     reg start_in_4_5;
     wire start_out_4_5;

     reg swap_in_4_5;
     wire swap_out_4_5;

     reg [1:0] op_in_4_5;
     wire [1:0] op_out_4_5;

     wire r_4_5;

     reg data_in_4_5;
     wire data_out_4_5;

     reg pivot_in_4_5;
     wire pivot_out_4_5;

     always @(posedge clk) begin
         op_in_4_5 <= op_out_4_4;
         pivot_in_4_5 <= pivot_out_4_4;
         start_in_4_5 <= start_out_4_4;
         swap_in_4_5 <= swap_out_4_4;
     end

     always @(posedge clk) begin
         data_in_4_5 <= data_out_3_5;
     end
  
     processor_AB AB_4_5 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_5),
       .start_in   (start_in_4_5),
       .swap_in   (swap_in_4_5),
       .op_in      (op_in_4_5),
       .pivot_in   (pivot_in_4_5),
       .start_out  (start_out_4_5),
       .swap_out   (swap_out_4_5),
       .data_out   (data_out_4_5),
       .op_out     (op_out_4_5),
       .pivot_out  (pivot_out_4_5),
       .r          (r_4_5)
     );

  // row 4, col 6

     reg start_in_4_6;
     wire start_out_4_6;

     reg swap_in_4_6;
     wire swap_out_4_6;

     reg [1:0] op_in_4_6;
     wire [1:0] op_out_4_6;

     wire r_4_6;

     reg data_in_4_6;
     wire data_out_4_6;

     reg pivot_in_4_6;
     wire pivot_out_4_6;

     always @(posedge clk) begin
         op_in_4_6 <= op_out_4_5;
         pivot_in_4_6 <= pivot_out_4_5;
         start_in_4_6 <= start_out_4_5;
         swap_in_4_6 <= swap_out_4_5;
     end

     always @(posedge clk) begin
         data_in_4_6 <= data_out_3_6;
     end
  
     processor_AB AB_4_6 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_6),
       .start_in   (start_in_4_6),
       .swap_in   (swap_in_4_6),
       .op_in      (op_in_4_6),
       .pivot_in   (pivot_in_4_6),
       .start_out  (start_out_4_6),
       .swap_out   (swap_out_4_6),
       .data_out   (data_out_4_6),
       .op_out     (op_out_4_6),
       .pivot_out  (pivot_out_4_6),
       .r          (r_4_6)
     );

  // row 4, col 7

     reg start_in_4_7;
     wire start_out_4_7;

     reg swap_in_4_7;
     wire swap_out_4_7;

     reg [1:0] op_in_4_7;
     wire [1:0] op_out_4_7;

     wire r_4_7;

     reg data_in_4_7;
     wire data_out_4_7;

     reg pivot_in_4_7;
     wire pivot_out_4_7;

     always @(posedge clk) begin
         op_in_4_7 <= op_out_4_6;
         pivot_in_4_7 <= pivot_out_4_6;
         start_in_4_7 <= start_out_4_6;
         swap_in_4_7 <= swap_out_4_6;
     end

     always @(posedge clk) begin
         data_in_4_7 <= data_out_3_7;
     end
  
     processor_AB AB_4_7 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_7),
       .start_in   (start_in_4_7),
       .swap_in   (swap_in_4_7),
       .op_in      (op_in_4_7),
       .pivot_in   (pivot_in_4_7),
       .start_out  (start_out_4_7),
       .swap_out   (swap_out_4_7),
       .data_out   (data_out_4_7),
       .op_out     (op_out_4_7),
       .pivot_out  (pivot_out_4_7),
       .r          (r_4_7)
     );

  // row 4, col 8

     reg start_in_4_8;
     wire start_out_4_8;

     reg swap_in_4_8;
     wire swap_out_4_8;

     reg [1:0] op_in_4_8;
     wire [1:0] op_out_4_8;

     wire r_4_8;

     reg data_in_4_8;
     wire data_out_4_8;

     reg pivot_in_4_8;
     wire pivot_out_4_8;

     always @(posedge clk) begin
         op_in_4_8 <= op_out_4_7;
         pivot_in_4_8 <= pivot_out_4_7;
         start_in_4_8 <= start_out_4_7;
         swap_in_4_8 <= swap_out_4_7;
     end

     always @(posedge clk) begin
         data_in_4_8 <= data_out_3_8;
     end
  
     processor_AB AB_4_8 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_8),
       .start_in   (start_in_4_8),
       .swap_in   (swap_in_4_8),
       .op_in      (op_in_4_8),
       .pivot_in   (pivot_in_4_8),
       .start_out  (start_out_4_8),
       .swap_out   (swap_out_4_8),
       .data_out   (data_out_4_8),
       .op_out     (op_out_4_8),
       .pivot_out  (pivot_out_4_8),
       .r          (r_4_8)
     );

  // row 4, col 9

     reg start_in_4_9;
     wire start_out_4_9;

     reg swap_in_4_9;
     wire swap_out_4_9;

     reg [1:0] op_in_4_9;
     wire [1:0] op_out_4_9;

     wire r_4_9;

     reg data_in_4_9;
     wire data_out_4_9;

     reg pivot_in_4_9;
     wire pivot_out_4_9;

     always @(posedge clk) begin
         op_in_4_9 <= op_out_4_8;
         pivot_in_4_9 <= pivot_out_4_8;
         start_in_4_9 <= start_out_4_8;
         swap_in_4_9 <= swap_out_4_8;
     end

     always @(posedge clk) begin
         data_in_4_9 <= data_out_3_9;
     end
  
     processor_AB AB_4_9 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_9),
       .start_in   (start_in_4_9),
       .swap_in   (swap_in_4_9),
       .op_in      (op_in_4_9),
       .pivot_in   (pivot_in_4_9),
       .start_out  (start_out_4_9),
       .swap_out   (swap_out_4_9),
       .data_out   (data_out_4_9),
       .op_out     (op_out_4_9),
       .pivot_out  (pivot_out_4_9),
       .r          (r_4_9)
     );

  // row 4, col 10

     reg start_in_4_10;
     wire start_out_4_10;

     reg swap_in_4_10;
     wire swap_out_4_10;

     reg [1:0] op_in_4_10;
     wire [1:0] op_out_4_10;

     wire r_4_10;

     reg data_in_4_10;
     wire data_out_4_10;

     reg pivot_in_4_10;
     wire pivot_out_4_10;

     always @(posedge clk) begin
         op_in_4_10 <= op_out_4_9;
         pivot_in_4_10 <= pivot_out_4_9;
         start_in_4_10 <= start_out_4_9;
         swap_in_4_10 <= swap_out_4_9;
     end

     always @(posedge clk) begin
         data_in_4_10 <= data_out_3_10;
     end
  
     processor_AB AB_4_10 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_10),
       .start_in   (start_in_4_10),
       .swap_in   (swap_in_4_10),
       .op_in      (op_in_4_10),
       .pivot_in   (pivot_in_4_10),
       .start_out  (start_out_4_10),
       .swap_out   (swap_out_4_10),
       .data_out   (data_out_4_10),
       .op_out     (op_out_4_10),
       .pivot_out  (pivot_out_4_10),
       .r          (r_4_10)
     );

  // row 4, col 11

     reg start_in_4_11;
     wire start_out_4_11;

     reg swap_in_4_11;
     wire swap_out_4_11;

     reg [1:0] op_in_4_11;
     wire [1:0] op_out_4_11;

     wire r_4_11;

     reg data_in_4_11;
     wire data_out_4_11;

     reg pivot_in_4_11;
     wire pivot_out_4_11;

     always @(posedge clk) begin
         op_in_4_11 <= op_out_4_10;
         pivot_in_4_11 <= pivot_out_4_10;
         start_in_4_11 <= start_out_4_10;
         swap_in_4_11 <= swap_out_4_10;
     end

     always @(posedge clk) begin
         data_in_4_11 <= data_out_3_11;
     end
  
     processor_AB AB_4_11 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_11),
       .start_in   (start_in_4_11),
       .swap_in   (swap_in_4_11),
       .op_in      (op_in_4_11),
       .pivot_in   (pivot_in_4_11),
       .start_out  (start_out_4_11),
       .swap_out   (swap_out_4_11),
       .data_out   (data_out_4_11),
       .op_out     (op_out_4_11),
       .pivot_out  (pivot_out_4_11),
       .r          (r_4_11)
     );

  // row 4, col 12

     reg start_in_4_12;
     wire start_out_4_12;

     reg swap_in_4_12;
     wire swap_out_4_12;

     reg [1:0] op_in_4_12;
     wire [1:0] op_out_4_12;

     wire r_4_12;

     reg data_in_4_12;
     wire data_out_4_12;

     reg pivot_in_4_12;
     wire pivot_out_4_12;

     always @(posedge clk) begin
         op_in_4_12 <= op_out_4_11;
         pivot_in_4_12 <= pivot_out_4_11;
         start_in_4_12 <= start_out_4_11;
         swap_in_4_12 <= swap_out_4_11;
     end

     always @(posedge clk) begin
         data_in_4_12 <= data_out_3_12;
     end
  
     processor_AB AB_4_12 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_12),
       .start_in   (start_in_4_12),
       .swap_in   (swap_in_4_12),
       .op_in      (op_in_4_12),
       .pivot_in   (pivot_in_4_12),
       .start_out  (start_out_4_12),
       .swap_out   (swap_out_4_12),
       .data_out   (data_out_4_12),
       .op_out     (op_out_4_12),
       .pivot_out  (pivot_out_4_12),
       .r          (r_4_12)
     );

  // row 4, col 13

     reg start_in_4_13;
     wire start_out_4_13;

     reg swap_in_4_13;
     wire swap_out_4_13;

     reg [1:0] op_in_4_13;
     wire [1:0] op_out_4_13;

     wire r_4_13;

     reg data_in_4_13;
     wire data_out_4_13;

     reg pivot_in_4_13;
     wire pivot_out_4_13;

     always @(posedge clk) begin
         op_in_4_13 <= op_out_4_12;
         pivot_in_4_13 <= pivot_out_4_12;
         start_in_4_13 <= start_out_4_12;
         swap_in_4_13 <= swap_out_4_12;
     end

     always @(posedge clk) begin
         data_in_4_13 <= data_out_3_13;
     end
  
     processor_AB AB_4_13 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_13),
       .start_in   (start_in_4_13),
       .swap_in   (swap_in_4_13),
       .op_in      (op_in_4_13),
       .pivot_in   (pivot_in_4_13),
       .start_out  (start_out_4_13),
       .swap_out   (swap_out_4_13),
       .data_out   (data_out_4_13),
       .op_out     (op_out_4_13),
       .pivot_out  (pivot_out_4_13),
       .r          (r_4_13)
     );

  // row 4, col 14

     reg start_in_4_14;
     wire start_out_4_14;

     reg swap_in_4_14;
     wire swap_out_4_14;

     reg [1:0] op_in_4_14;
     wire [1:0] op_out_4_14;

     wire r_4_14;

     reg data_in_4_14;
     wire data_out_4_14;

     reg pivot_in_4_14;
     wire pivot_out_4_14;

     always @(posedge clk) begin
         op_in_4_14 <= op_out_4_13;
         pivot_in_4_14 <= pivot_out_4_13;
         start_in_4_14 <= start_out_4_13;
         swap_in_4_14 <= swap_out_4_13;
     end

     always @(posedge clk) begin
         data_in_4_14 <= data_out_3_14;
     end
  
     processor_AB AB_4_14 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_14),
       .start_in   (start_in_4_14),
       .swap_in   (swap_in_4_14),
       .op_in      (op_in_4_14),
       .pivot_in   (pivot_in_4_14),
       .start_out  (start_out_4_14),
       .swap_out   (swap_out_4_14),
       .data_out   (data_out_4_14),
       .op_out     (op_out_4_14),
       .pivot_out  (pivot_out_4_14),
       .r          (r_4_14)
     );

  // row 4, col 15

     reg start_in_4_15;
     wire start_out_4_15;

     reg swap_in_4_15;
     wire swap_out_4_15;

     reg [1:0] op_in_4_15;
     wire [1:0] op_out_4_15;

     wire r_4_15;

     reg data_in_4_15;
     wire data_out_4_15;

     reg pivot_in_4_15;
     wire pivot_out_4_15;

     always @(posedge clk) begin
         op_in_4_15 <= op_out_4_14;
         pivot_in_4_15 <= pivot_out_4_14;
         start_in_4_15 <= start_out_4_14;
         swap_in_4_15 <= swap_out_4_14;
     end

     always @(posedge clk) begin
         data_in_4_15 <= data_out_3_15;
     end
  
     processor_AB AB_4_15 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_15),
       .start_in   (start_in_4_15),
       .swap_in   (swap_in_4_15),
       .op_in      (op_in_4_15),
       .pivot_in   (pivot_in_4_15),
       .start_out  (start_out_4_15),
       .swap_out   (swap_out_4_15),
       .data_out   (data_out_4_15),
       .op_out     (op_out_4_15),
       .pivot_out  (pivot_out_4_15),
       .r          (r_4_15)
     );

  // row 4, col 16

     reg start_in_4_16;
     wire start_out_4_16;

     reg swap_in_4_16;
     wire swap_out_4_16;

     reg [1:0] op_in_4_16;
     wire [1:0] op_out_4_16;

     wire r_4_16;

     reg data_in_4_16;
     wire data_out_4_16;

     reg pivot_in_4_16;
     wire pivot_out_4_16;

     always @(posedge clk) begin
         op_in_4_16 <= op_out_4_15;
         pivot_in_4_16 <= pivot_out_4_15;
         start_in_4_16 <= start_out_4_15;
         swap_in_4_16 <= swap_out_4_15;
     end

     always @(posedge clk) begin
         data_in_4_16 <= data_out_3_16;
     end
  
     processor_AB AB_4_16 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_16),
       .start_in   (start_in_4_16),
       .swap_in   (swap_in_4_16),
       .op_in      (op_in_4_16),
       .pivot_in   (pivot_in_4_16),
       .start_out  (start_out_4_16),
       .swap_out   (swap_out_4_16),
       .data_out   (data_out_4_16),
       .op_out     (op_out_4_16),
       .pivot_out  (pivot_out_4_16),
       .r          (r_4_16)
     );

  // row 4, col 17

     reg start_in_4_17;
     wire start_out_4_17;

     reg swap_in_4_17;
     wire swap_out_4_17;

     reg [1:0] op_in_4_17;
     wire [1:0] op_out_4_17;

     wire r_4_17;

     reg data_in_4_17;
     wire data_out_4_17;

     reg pivot_in_4_17;
     wire pivot_out_4_17;

     always @(posedge clk) begin
         op_in_4_17 <= op_out_4_16;
         pivot_in_4_17 <= pivot_out_4_16;
         start_in_4_17 <= start_out_4_16;
         swap_in_4_17 <= swap_out_4_16;
     end

     always @(posedge clk) begin
         data_in_4_17 <= data_out_3_17;
     end
  
     processor_AB AB_4_17 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_17),
       .start_in   (start_in_4_17),
       .swap_in   (swap_in_4_17),
       .op_in      (op_in_4_17),
       .pivot_in   (pivot_in_4_17),
       .start_out  (start_out_4_17),
       .swap_out   (swap_out_4_17),
       .data_out   (data_out_4_17),
       .op_out     (op_out_4_17),
       .pivot_out  (pivot_out_4_17),
       .r          (r_4_17)
     );

  // row 4, col 18

     reg start_in_4_18;
     wire start_out_4_18;

     reg swap_in_4_18;
     wire swap_out_4_18;

     reg [1:0] op_in_4_18;
     wire [1:0] op_out_4_18;

     wire r_4_18;

     reg data_in_4_18;
     wire data_out_4_18;

     reg pivot_in_4_18;
     wire pivot_out_4_18;

     always @(posedge clk) begin
         op_in_4_18 <= op_out_4_17;
         pivot_in_4_18 <= pivot_out_4_17;
         start_in_4_18 <= start_out_4_17;
         swap_in_4_18 <= swap_out_4_17;
     end

     always @(posedge clk) begin
         data_in_4_18 <= data_out_3_18;
     end
  
     processor_AB AB_4_18 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_18),
       .start_in   (start_in_4_18),
       .swap_in   (swap_in_4_18),
       .op_in      (op_in_4_18),
       .pivot_in   (pivot_in_4_18),
       .start_out  (start_out_4_18),
       .swap_out   (swap_out_4_18),
       .data_out   (data_out_4_18),
       .op_out     (op_out_4_18),
       .pivot_out  (pivot_out_4_18),
       .r          (r_4_18)
     );

  // row 4, col 19

     reg start_in_4_19;
     wire start_out_4_19;

     reg swap_in_4_19;
     wire swap_out_4_19;

     reg [1:0] op_in_4_19;
     wire [1:0] op_out_4_19;

     wire r_4_19;

     reg data_in_4_19;
     wire data_out_4_19;

     reg pivot_in_4_19;
     wire pivot_out_4_19;

     always @(posedge clk) begin
         op_in_4_19 <= op_out_4_18;
         pivot_in_4_19 <= pivot_out_4_18;
         start_in_4_19 <= start_out_4_18;
         swap_in_4_19 <= swap_out_4_18;
     end

     always @(posedge clk) begin
         data_in_4_19 <= data_out_3_19;
     end
  
     processor_AB AB_4_19 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_19),
       .start_in   (start_in_4_19),
       .swap_in   (swap_in_4_19),
       .op_in      (op_in_4_19),
       .pivot_in   (pivot_in_4_19),
       .start_out  (start_out_4_19),
       .swap_out   (swap_out_4_19),
       .data_out   (data_out_4_19),
       .op_out     (op_out_4_19),
       .pivot_out  (pivot_out_4_19),
       .r          (r_4_19)
     );

  // row 4, col 20

     reg start_in_4_20;
     wire start_out_4_20;

     reg swap_in_4_20;
     wire swap_out_4_20;

     reg [1:0] op_in_4_20;
     wire [1:0] op_out_4_20;

     wire r_4_20;

     reg data_in_4_20;
     wire data_out_4_20;

     reg pivot_in_4_20;
     wire pivot_out_4_20;

     always @(posedge clk) begin
         op_in_4_20 <= op_out_4_19;
         pivot_in_4_20 <= pivot_out_4_19;
         start_in_4_20 <= start_out_4_19;
         swap_in_4_20 <= swap_out_4_19;
     end

     always @(posedge clk) begin
         data_in_4_20 <= data_out_3_20;
     end
  
     processor_AB AB_4_20 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_20),
       .start_in   (start_in_4_20),
       .swap_in   (swap_in_4_20),
       .op_in      (op_in_4_20),
       .pivot_in   (pivot_in_4_20),
       .start_out  (start_out_4_20),
       .swap_out   (swap_out_4_20),
       .data_out   (data_out_4_20),
       .op_out     (op_out_4_20),
       .pivot_out  (pivot_out_4_20),
       .r          (r_4_20)
     );

  // row 4, col 21

     reg start_in_4_21;
     wire start_out_4_21;

     reg swap_in_4_21;
     wire swap_out_4_21;

     reg [1:0] op_in_4_21;
     wire [1:0] op_out_4_21;

     wire r_4_21;

     reg data_in_4_21;
     wire data_out_4_21;

     reg pivot_in_4_21;
     wire pivot_out_4_21;

     always @(posedge clk) begin
         op_in_4_21 <= op_out_4_20;
         pivot_in_4_21 <= pivot_out_4_20;
         start_in_4_21 <= start_out_4_20;
         swap_in_4_21 <= swap_out_4_20;
     end

     always @(posedge clk) begin
         data_in_4_21 <= data_out_3_21;
     end
  
     processor_AB AB_4_21 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_21),
       .start_in   (start_in_4_21),
       .swap_in   (swap_in_4_21),
       .op_in      (op_in_4_21),
       .pivot_in   (pivot_in_4_21),
       .start_out  (start_out_4_21),
       .swap_out   (swap_out_4_21),
       .data_out   (data_out_4_21),
       .op_out     (op_out_4_21),
       .pivot_out  (pivot_out_4_21),
       .r          (r_4_21)
     );

  // row 4, col 22

     reg start_in_4_22;
     wire start_out_4_22;

     reg swap_in_4_22;
     wire swap_out_4_22;

     reg [1:0] op_in_4_22;
     wire [1:0] op_out_4_22;

     wire r_4_22;

     reg data_in_4_22;
     wire data_out_4_22;

     reg pivot_in_4_22;
     wire pivot_out_4_22;

     always @(posedge clk) begin
         op_in_4_22 <= op_out_4_21;
         pivot_in_4_22 <= pivot_out_4_21;
         start_in_4_22 <= start_out_4_21;
         swap_in_4_22 <= swap_out_4_21;
     end

     always @(posedge clk) begin
         data_in_4_22 <= data_out_3_22;
     end
  
     processor_AB AB_4_22 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_22),
       .start_in   (start_in_4_22),
       .swap_in   (swap_in_4_22),
       .op_in      (op_in_4_22),
       .pivot_in   (pivot_in_4_22),
       .start_out  (start_out_4_22),
       .swap_out   (swap_out_4_22),
       .data_out   (data_out_4_22),
       .op_out     (op_out_4_22),
       .pivot_out  (pivot_out_4_22),
       .r          (r_4_22)
     );

  // row 4, col 23

     reg start_in_4_23;
     wire start_out_4_23;

     reg swap_in_4_23;
     wire swap_out_4_23;

     reg [1:0] op_in_4_23;
     wire [1:0] op_out_4_23;

     wire r_4_23;

     reg data_in_4_23;
     wire data_out_4_23;

     reg pivot_in_4_23;
     wire pivot_out_4_23;

     always @(posedge clk) begin
         op_in_4_23 <= op_out_4_22;
         pivot_in_4_23 <= pivot_out_4_22;
         start_in_4_23 <= start_out_4_22;
         swap_in_4_23 <= swap_out_4_22;
     end

     always @(posedge clk) begin
         data_in_4_23 <= data_out_3_23;
     end
  
     processor_AB AB_4_23 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_23),
       .start_in   (start_in_4_23),
       .swap_in   (swap_in_4_23),
       .op_in      (op_in_4_23),
       .pivot_in   (pivot_in_4_23),
       .start_out  (start_out_4_23),
       .swap_out   (swap_out_4_23),
       .data_out   (data_out_4_23),
       .op_out     (op_out_4_23),
       .pivot_out  (pivot_out_4_23),
       .r          (r_4_23)
     );

  // row 4, col 24

     reg start_in_4_24;
     wire start_out_4_24;

     reg swap_in_4_24;
     wire swap_out_4_24;

     reg [1:0] op_in_4_24;
     wire [1:0] op_out_4_24;

     wire r_4_24;

     reg data_in_4_24;
     wire data_out_4_24;

     reg pivot_in_4_24;
     wire pivot_out_4_24;

     always @(posedge clk) begin
         op_in_4_24 <= op_out_4_23;
         pivot_in_4_24 <= pivot_out_4_23;
         start_in_4_24 <= start_out_4_23;
         swap_in_4_24 <= swap_out_4_23;
     end

     always @(posedge clk) begin
         data_in_4_24 <= data_out_3_24;
     end
  
     processor_AB AB_4_24 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_24),
       .start_in   (start_in_4_24),
       .swap_in   (swap_in_4_24),
       .op_in      (op_in_4_24),
       .pivot_in   (pivot_in_4_24),
       .start_out  (start_out_4_24),
       .swap_out   (swap_out_4_24),
       .data_out   (data_out_4_24),
       .op_out     (op_out_4_24),
       .pivot_out  (pivot_out_4_24),
       .r          (r_4_24)
     );

  // row 4, col 25

     reg start_in_4_25;
     wire start_out_4_25;

     reg swap_in_4_25;
     wire swap_out_4_25;

     reg [1:0] op_in_4_25;
     wire [1:0] op_out_4_25;

     wire r_4_25;

     reg data_in_4_25;
     wire data_out_4_25;

     reg pivot_in_4_25;
     wire pivot_out_4_25;

     always @(posedge clk) begin
         op_in_4_25 <= op_out_4_24;
         pivot_in_4_25 <= pivot_out_4_24;
         start_in_4_25 <= start_out_4_24;
         swap_in_4_25 <= swap_out_4_24;
     end

     always @(posedge clk) begin
         data_in_4_25 <= data_out_3_25;
     end
  
     processor_AB AB_4_25 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_25),
       .start_in   (start_in_4_25),
       .swap_in   (swap_in_4_25),
       .op_in      (op_in_4_25),
       .pivot_in   (pivot_in_4_25),
       .start_out  (start_out_4_25),
       .swap_out   (swap_out_4_25),
       .data_out   (data_out_4_25),
       .op_out     (op_out_4_25),
       .pivot_out  (pivot_out_4_25),
       .r          (r_4_25)
     );

  // row 4, col 26

     reg start_in_4_26;
     wire start_out_4_26;

     reg swap_in_4_26;
     wire swap_out_4_26;

     reg [1:0] op_in_4_26;
     wire [1:0] op_out_4_26;

     wire r_4_26;

     reg data_in_4_26;
     wire data_out_4_26;

     reg pivot_in_4_26;
     wire pivot_out_4_26;

     always @(posedge clk) begin
         op_in_4_26 <= op_out_4_25;
         pivot_in_4_26 <= pivot_out_4_25;
         start_in_4_26 <= start_out_4_25;
         swap_in_4_26 <= swap_out_4_25;
     end

     always @(posedge clk) begin
         data_in_4_26 <= data_out_3_26;
     end
  
     processor_AB AB_4_26 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_26),
       .start_in   (start_in_4_26),
       .swap_in   (swap_in_4_26),
       .op_in      (op_in_4_26),
       .pivot_in   (pivot_in_4_26),
       .start_out  (start_out_4_26),
       .swap_out   (swap_out_4_26),
       .data_out   (data_out_4_26),
       .op_out     (op_out_4_26),
       .pivot_out  (pivot_out_4_26),
       .r          (r_4_26)
     );

  // row 4, col 27

     reg start_in_4_27;
     wire start_out_4_27;

     reg swap_in_4_27;
     wire swap_out_4_27;

     reg [1:0] op_in_4_27;
     wire [1:0] op_out_4_27;

     wire r_4_27;

     reg data_in_4_27;
     wire data_out_4_27;

     reg pivot_in_4_27;
     wire pivot_out_4_27;

     always @(posedge clk) begin
         op_in_4_27 <= op_out_4_26;
         pivot_in_4_27 <= pivot_out_4_26;
         start_in_4_27 <= start_out_4_26;
         swap_in_4_27 <= swap_out_4_26;
     end

     always @(posedge clk) begin
         data_in_4_27 <= data_out_3_27;
     end
  
     processor_AB AB_4_27 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_27),
       .start_in   (start_in_4_27),
       .swap_in   (swap_in_4_27),
       .op_in      (op_in_4_27),
       .pivot_in   (pivot_in_4_27),
       .start_out  (start_out_4_27),
       .swap_out   (swap_out_4_27),
       .data_out   (data_out_4_27),
       .op_out     (op_out_4_27),
       .pivot_out  (pivot_out_4_27),
       .r          (r_4_27)
     );

  // row 4, col 28

     reg start_in_4_28;
     wire start_out_4_28;

     reg swap_in_4_28;
     wire swap_out_4_28;

     reg [1:0] op_in_4_28;
     wire [1:0] op_out_4_28;

     wire r_4_28;

     reg data_in_4_28;
     wire data_out_4_28;

     reg pivot_in_4_28;
     wire pivot_out_4_28;

     always @(posedge clk) begin
         op_in_4_28 <= op_out_4_27;
         pivot_in_4_28 <= pivot_out_4_27;
         start_in_4_28 <= start_out_4_27;
         swap_in_4_28 <= swap_out_4_27;
     end

     always @(posedge clk) begin
         data_in_4_28 <= data_out_3_28;
     end
  
     processor_AB AB_4_28 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_28),
       .start_in   (start_in_4_28),
       .swap_in   (swap_in_4_28),
       .op_in      (op_in_4_28),
       .pivot_in   (pivot_in_4_28),
       .start_out  (start_out_4_28),
       .swap_out   (swap_out_4_28),
       .data_out   (data_out_4_28),
       .op_out     (op_out_4_28),
       .pivot_out  (pivot_out_4_28),
       .r          (r_4_28)
     );

  // row 4, col 29

     reg start_in_4_29;
     wire start_out_4_29;

     reg swap_in_4_29;
     wire swap_out_4_29;

     reg [1:0] op_in_4_29;
     wire [1:0] op_out_4_29;

     wire r_4_29;

     reg data_in_4_29;
     wire data_out_4_29;

     reg pivot_in_4_29;
     wire pivot_out_4_29;

     always @(posedge clk) begin
         op_in_4_29 <= op_out_4_28;
         pivot_in_4_29 <= pivot_out_4_28;
         start_in_4_29 <= start_out_4_28;
         swap_in_4_29 <= swap_out_4_28;
     end

     always @(posedge clk) begin
         data_in_4_29 <= data_out_3_29;
     end
  
     processor_AB AB_4_29 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_29),
       .start_in   (start_in_4_29),
       .swap_in   (swap_in_4_29),
       .op_in      (op_in_4_29),
       .pivot_in   (pivot_in_4_29),
       .start_out  (start_out_4_29),
       .swap_out   (swap_out_4_29),
       .data_out   (data_out_4_29),
       .op_out     (op_out_4_29),
       .pivot_out  (pivot_out_4_29),
       .r          (r_4_29)
     );

  // row 4, col 30

     reg start_in_4_30;
     wire start_out_4_30;

     reg swap_in_4_30;
     wire swap_out_4_30;

     reg [1:0] op_in_4_30;
     wire [1:0] op_out_4_30;

     wire r_4_30;

     reg data_in_4_30;
     wire data_out_4_30;

     reg pivot_in_4_30;
     wire pivot_out_4_30;

     always @(posedge clk) begin
         op_in_4_30 <= op_out_4_29;
         pivot_in_4_30 <= pivot_out_4_29;
         start_in_4_30 <= start_out_4_29;
         swap_in_4_30 <= swap_out_4_29;
     end

     always @(posedge clk) begin
         data_in_4_30 <= data_out_3_30;
     end
  
     processor_AB AB_4_30 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_30),
       .start_in   (start_in_4_30),
       .swap_in   (swap_in_4_30),
       .op_in      (op_in_4_30),
       .pivot_in   (pivot_in_4_30),
       .start_out  (start_out_4_30),
       .swap_out   (swap_out_4_30),
       .data_out   (data_out_4_30),
       .op_out     (op_out_4_30),
       .pivot_out  (pivot_out_4_30),
       .r          (r_4_30)
     );

  // row 4, col 31

     reg start_in_4_31;
     wire start_out_4_31;

     reg swap_in_4_31;
     wire swap_out_4_31;

     reg [1:0] op_in_4_31;
     wire [1:0] op_out_4_31;

     wire r_4_31;

     reg data_in_4_31;
     wire data_out_4_31;

     reg pivot_in_4_31;
     wire pivot_out_4_31;

     always @(posedge clk) begin
         op_in_4_31 <= op_out_4_30;
         pivot_in_4_31 <= pivot_out_4_30;
         start_in_4_31 <= start_out_4_30;
         swap_in_4_31 <= swap_out_4_30;
     end

     always @(posedge clk) begin
         data_in_4_31 <= data_out_3_31;
     end
  
     processor_AB AB_4_31 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_31),
       .start_in   (start_in_4_31),
       .swap_in   (swap_in_4_31),
       .op_in      (op_in_4_31),
       .pivot_in   (pivot_in_4_31),
       .start_out  (start_out_4_31),
       .swap_out   (swap_out_4_31),
       .data_out   (data_out_4_31),
       .op_out     (op_out_4_31),
       .pivot_out  (pivot_out_4_31),
       .r          (r_4_31)
     );

  // row 4, col 32

     reg start_in_4_32;
     wire start_out_4_32;

     reg swap_in_4_32;
     wire swap_out_4_32;

     reg [1:0] op_in_4_32;
     wire [1:0] op_out_4_32;

     wire r_4_32;

     reg data_in_4_32;
     wire data_out_4_32;

     reg pivot_in_4_32;
     wire pivot_out_4_32;

     always @(posedge clk) begin
         op_in_4_32 <= op_out_4_31;
         pivot_in_4_32 <= pivot_out_4_31;
         start_in_4_32 <= start_out_4_31;
         swap_in_4_32 <= swap_out_4_31;
     end

     always @(posedge clk) begin
         data_in_4_32 <= data_out_3_32;
     end
  
     processor_AB AB_4_32 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_32),
       .start_in   (start_in_4_32),
       .swap_in   (swap_in_4_32),
       .op_in      (op_in_4_32),
       .pivot_in   (pivot_in_4_32),
       .start_out  (start_out_4_32),
       .swap_out   (swap_out_4_32),
       .data_out   (data_out_4_32),
       .op_out     (op_out_4_32),
       .pivot_out  (pivot_out_4_32),
       .r          (r_4_32)
     );

  // row 4, col 33

     reg start_in_4_33;
     wire start_out_4_33;

     reg swap_in_4_33;
     wire swap_out_4_33;

     reg [1:0] op_in_4_33;
     wire [1:0] op_out_4_33;

     wire r_4_33;

     reg data_in_4_33;
     wire data_out_4_33;

     reg pivot_in_4_33;
     wire pivot_out_4_33;

     always @(posedge clk) begin
         op_in_4_33 <= op_out_4_32;
         pivot_in_4_33 <= pivot_out_4_32;
         start_in_4_33 <= start_out_4_32;
         swap_in_4_33 <= swap_out_4_32;
     end

     always @(posedge clk) begin
         data_in_4_33 <= data_out_3_33;
     end
  
     processor_AB AB_4_33 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_33),
       .start_in   (start_in_4_33),
       .swap_in   (swap_in_4_33),
       .op_in      (op_in_4_33),
       .pivot_in   (pivot_in_4_33),
       .start_out  (start_out_4_33),
       .swap_out   (swap_out_4_33),
       .data_out   (data_out_4_33),
       .op_out     (op_out_4_33),
       .pivot_out  (pivot_out_4_33),
       .r          (r_4_33)
     );

  // row 4, col 34

     reg start_in_4_34;
     wire start_out_4_34;

     reg swap_in_4_34;
     wire swap_out_4_34;

     reg [1:0] op_in_4_34;
     wire [1:0] op_out_4_34;

     wire r_4_34;

     reg data_in_4_34;
     wire data_out_4_34;

     reg pivot_in_4_34;
     wire pivot_out_4_34;

     always @(posedge clk) begin
         op_in_4_34 <= op_out_4_33;
         pivot_in_4_34 <= pivot_out_4_33;
         start_in_4_34 <= start_out_4_33;
         swap_in_4_34 <= swap_out_4_33;
     end

     always @(posedge clk) begin
         data_in_4_34 <= data_out_3_34;
     end
  
     processor_AB AB_4_34 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_34),
       .start_in   (start_in_4_34),
       .swap_in   (swap_in_4_34),
       .op_in      (op_in_4_34),
       .pivot_in   (pivot_in_4_34),
       .start_out  (start_out_4_34),
       .swap_out   (swap_out_4_34),
       .data_out   (data_out_4_34),
       .op_out     (op_out_4_34),
       .pivot_out  (pivot_out_4_34),
       .r          (r_4_34)
     );

  // row 4, col 35

     reg start_in_4_35;
     wire start_out_4_35;

     reg swap_in_4_35;
     wire swap_out_4_35;

     reg [1:0] op_in_4_35;
     wire [1:0] op_out_4_35;

     wire r_4_35;

     reg data_in_4_35;
     wire data_out_4_35;

     reg pivot_in_4_35;
     wire pivot_out_4_35;

     always @(posedge clk) begin
         op_in_4_35 <= op_out_4_34;
         pivot_in_4_35 <= pivot_out_4_34;
         start_in_4_35 <= start_out_4_34;
         swap_in_4_35 <= swap_out_4_34;
     end

     always @(posedge clk) begin
         data_in_4_35 <= data_out_3_35;
     end
  
     processor_AB AB_4_35 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_35),
       .start_in   (start_in_4_35),
       .swap_in   (swap_in_4_35),
       .op_in      (op_in_4_35),
       .pivot_in   (pivot_in_4_35),
       .start_out  (start_out_4_35),
       .swap_out   (swap_out_4_35),
       .data_out   (data_out_4_35),
       .op_out     (op_out_4_35),
       .pivot_out  (pivot_out_4_35),
       .r          (r_4_35)
     );

  // row 4, col 36

     reg start_in_4_36;
     wire start_out_4_36;

     reg swap_in_4_36;
     wire swap_out_4_36;

     reg [1:0] op_in_4_36;
     wire [1:0] op_out_4_36;

     wire r_4_36;

     reg data_in_4_36;
     wire data_out_4_36;

     reg pivot_in_4_36;
     wire pivot_out_4_36;

     always @(posedge clk) begin
         op_in_4_36 <= op_out_4_35;
         pivot_in_4_36 <= pivot_out_4_35;
         start_in_4_36 <= start_out_4_35;
         swap_in_4_36 <= swap_out_4_35;
     end

     always @(posedge clk) begin
         data_in_4_36 <= data_out_3_36;
     end
  
     processor_AB AB_4_36 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_36),
       .start_in   (start_in_4_36),
       .swap_in   (swap_in_4_36),
       .op_in      (op_in_4_36),
       .pivot_in   (pivot_in_4_36),
       .start_out  (start_out_4_36),
       .swap_out   (swap_out_4_36),
       .data_out   (data_out_4_36),
       .op_out     (op_out_4_36),
       .pivot_out  (pivot_out_4_36),
       .r          (r_4_36)
     );

  // row 4, col 37

     reg start_in_4_37;
     wire start_out_4_37;

     reg swap_in_4_37;
     wire swap_out_4_37;

     reg [1:0] op_in_4_37;
     wire [1:0] op_out_4_37;

     wire r_4_37;

     reg data_in_4_37;
     wire data_out_4_37;

     reg pivot_in_4_37;
     wire pivot_out_4_37;

     always @(posedge clk) begin
         op_in_4_37 <= op_out_4_36;
         pivot_in_4_37 <= pivot_out_4_36;
         start_in_4_37 <= start_out_4_36;
         swap_in_4_37 <= swap_out_4_36;
     end

     always @(posedge clk) begin
         data_in_4_37 <= data_out_3_37;
     end
  
     processor_AB AB_4_37 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_37),
       .start_in   (start_in_4_37),
       .swap_in   (swap_in_4_37),
       .op_in      (op_in_4_37),
       .pivot_in   (pivot_in_4_37),
       .start_out  (start_out_4_37),
       .swap_out   (swap_out_4_37),
       .data_out   (data_out_4_37),
       .op_out     (op_out_4_37),
       .pivot_out  (pivot_out_4_37),
       .r          (r_4_37)
     );

  // row 4, col 38

     reg start_in_4_38;
     wire start_out_4_38;

     reg swap_in_4_38;
     wire swap_out_4_38;

     reg [1:0] op_in_4_38;
     wire [1:0] op_out_4_38;

     wire r_4_38;

     reg data_in_4_38;
     wire data_out_4_38;

     reg pivot_in_4_38;
     wire pivot_out_4_38;

     always @(posedge clk) begin
         op_in_4_38 <= op_out_4_37;
         pivot_in_4_38 <= pivot_out_4_37;
         start_in_4_38 <= start_out_4_37;
         swap_in_4_38 <= swap_out_4_37;
     end

     always @(posedge clk) begin
         data_in_4_38 <= data_out_3_38;
     end
  
     processor_AB AB_4_38 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_38),
       .start_in   (start_in_4_38),
       .swap_in   (swap_in_4_38),
       .op_in      (op_in_4_38),
       .pivot_in   (pivot_in_4_38),
       .start_out  (start_out_4_38),
       .swap_out   (swap_out_4_38),
       .data_out   (data_out_4_38),
       .op_out     (op_out_4_38),
       .pivot_out  (pivot_out_4_38),
       .r          (r_4_38)
     );

  // row 4, col 39

     reg start_in_4_39;
     wire start_out_4_39;

     reg swap_in_4_39;
     wire swap_out_4_39;

     reg [1:0] op_in_4_39;
     wire [1:0] op_out_4_39;

     wire r_4_39;

     reg data_in_4_39;
     wire data_out_4_39;

     reg pivot_in_4_39;
     wire pivot_out_4_39;

     always @(posedge clk) begin
         op_in_4_39 <= op_out_4_38;
         pivot_in_4_39 <= pivot_out_4_38;
         start_in_4_39 <= start_out_4_38;
         swap_in_4_39 <= swap_out_4_38;
     end

     always @(posedge clk) begin
         data_in_4_39 <= data_out_3_39;
     end
  
     processor_AB AB_4_39 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_39),
       .start_in   (start_in_4_39),
       .swap_in   (swap_in_4_39),
       .op_in      (op_in_4_39),
       .pivot_in   (pivot_in_4_39),
       .start_out  (start_out_4_39),
       .swap_out   (swap_out_4_39),
       .data_out   (data_out_4_39),
       .op_out     (op_out_4_39),
       .pivot_out  (pivot_out_4_39),
       .r          (r_4_39)
     );

  // row 4, col 40

     reg start_in_4_40;
     wire start_out_4_40;

     reg swap_in_4_40;
     wire swap_out_4_40;

     reg [1:0] op_in_4_40;
     wire [1:0] op_out_4_40;

     wire r_4_40;

     reg data_in_4_40;
     wire data_out_4_40;

     reg pivot_in_4_40;
     wire pivot_out_4_40;

     always @(posedge clk) begin
         op_in_4_40 <= op_out_4_39;
         pivot_in_4_40 <= pivot_out_4_39;
         start_in_4_40 <= start_out_4_39;
         swap_in_4_40 <= swap_out_4_39;
     end

     always @(posedge clk) begin
         data_in_4_40 <= data_out_3_40;
     end
  
     processor_AB AB_4_40 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_40),
       .start_in   (start_in_4_40),
       .swap_in   (swap_in_4_40),
       .op_in      (op_in_4_40),
       .pivot_in   (pivot_in_4_40),
       .start_out  (start_out_4_40),
       .swap_out   (swap_out_4_40),
       .data_out   (data_out_4_40),
       .op_out     (op_out_4_40),
       .pivot_out  (pivot_out_4_40),
       .r          (r_4_40)
     );

  // row 4, col 41

     reg start_in_4_41;
     wire start_out_4_41;

     reg swap_in_4_41;
     wire swap_out_4_41;

     reg [1:0] op_in_4_41;
     wire [1:0] op_out_4_41;

     wire r_4_41;

     reg data_in_4_41;
     wire data_out_4_41;

     reg pivot_in_4_41;
     wire pivot_out_4_41;

     always @(posedge clk) begin
         op_in_4_41 <= op_out_4_40;
         pivot_in_4_41 <= pivot_out_4_40;
         start_in_4_41 <= start_out_4_40;
         swap_in_4_41 <= swap_out_4_40;
     end

     always @(posedge clk) begin
         data_in_4_41 <= data_out_3_41;
     end
  
     processor_AB AB_4_41 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_41),
       .start_in   (start_in_4_41),
       .swap_in   (swap_in_4_41),
       .op_in      (op_in_4_41),
       .pivot_in   (pivot_in_4_41),
       .start_out  (start_out_4_41),
       .swap_out   (swap_out_4_41),
       .data_out   (data_out_4_41),
       .op_out     (op_out_4_41),
       .pivot_out  (pivot_out_4_41),
       .r          (r_4_41)
     );

  // row 4, col 42

     reg start_in_4_42;
     wire start_out_4_42;

     reg swap_in_4_42;
     wire swap_out_4_42;

     reg [1:0] op_in_4_42;
     wire [1:0] op_out_4_42;

     wire r_4_42;

     reg data_in_4_42;
     wire data_out_4_42;

     reg pivot_in_4_42;
     wire pivot_out_4_42;

     always @(posedge clk) begin
         op_in_4_42 <= op_out_4_41;
         pivot_in_4_42 <= pivot_out_4_41;
         start_in_4_42 <= start_out_4_41;
         swap_in_4_42 <= swap_out_4_41;
     end

     always @(posedge clk) begin
         data_in_4_42 <= data_out_3_42;
     end
  
     processor_AB AB_4_42 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_42),
       .start_in   (start_in_4_42),
       .swap_in   (swap_in_4_42),
       .op_in      (op_in_4_42),
       .pivot_in   (pivot_in_4_42),
       .start_out  (start_out_4_42),
       .swap_out   (swap_out_4_42),
       .data_out   (data_out_4_42),
       .op_out     (op_out_4_42),
       .pivot_out  (pivot_out_4_42),
       .r          (r_4_42)
     );

  // row 4, col 43

     reg start_in_4_43;
     wire start_out_4_43;

     reg swap_in_4_43;
     wire swap_out_4_43;

     reg [1:0] op_in_4_43;
     wire [1:0] op_out_4_43;

     wire r_4_43;

     reg data_in_4_43;
     wire data_out_4_43;

     reg pivot_in_4_43;
     wire pivot_out_4_43;

     always @(posedge clk) begin
         op_in_4_43 <= op_out_4_42;
         pivot_in_4_43 <= pivot_out_4_42;
         start_in_4_43 <= start_out_4_42;
         swap_in_4_43 <= swap_out_4_42;
     end

     always @(posedge clk) begin
         data_in_4_43 <= data_out_3_43;
     end
  
     processor_AB AB_4_43 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_43),
       .start_in   (start_in_4_43),
       .swap_in   (swap_in_4_43),
       .op_in      (op_in_4_43),
       .pivot_in   (pivot_in_4_43),
       .start_out  (start_out_4_43),
       .swap_out   (swap_out_4_43),
       .data_out   (data_out_4_43),
       .op_out     (op_out_4_43),
       .pivot_out  (pivot_out_4_43),
       .r          (r_4_43)
     );

  // row 4, col 44

     reg start_in_4_44;
     wire start_out_4_44;

     reg swap_in_4_44;
     wire swap_out_4_44;

     reg [1:0] op_in_4_44;
     wire [1:0] op_out_4_44;

     wire r_4_44;

     reg data_in_4_44;
     wire data_out_4_44;

     reg pivot_in_4_44;
     wire pivot_out_4_44;

     always @(posedge clk) begin
         op_in_4_44 <= op_out_4_43;
         pivot_in_4_44 <= pivot_out_4_43;
         start_in_4_44 <= start_out_4_43;
         swap_in_4_44 <= swap_out_4_43;
     end

     always @(posedge clk) begin
         data_in_4_44 <= data_out_3_44;
     end
  
     processor_AB AB_4_44 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_44),
       .start_in   (start_in_4_44),
       .swap_in   (swap_in_4_44),
       .op_in      (op_in_4_44),
       .pivot_in   (pivot_in_4_44),
       .start_out  (start_out_4_44),
       .swap_out   (swap_out_4_44),
       .data_out   (data_out_4_44),
       .op_out     (op_out_4_44),
       .pivot_out  (pivot_out_4_44),
       .r          (r_4_44)
     );

  // row 4, col 45

     reg start_in_4_45;
     wire start_out_4_45;

     reg swap_in_4_45;
     wire swap_out_4_45;

     reg [1:0] op_in_4_45;
     wire [1:0] op_out_4_45;

     wire r_4_45;

     reg data_in_4_45;
     wire data_out_4_45;

     reg pivot_in_4_45;
     wire pivot_out_4_45;

     always @(posedge clk) begin
         op_in_4_45 <= op_out_4_44;
         pivot_in_4_45 <= pivot_out_4_44;
         start_in_4_45 <= start_out_4_44;
         swap_in_4_45 <= swap_out_4_44;
     end

     always @(posedge clk) begin
         data_in_4_45 <= data_out_3_45;
     end
  
     processor_AB AB_4_45 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_45),
       .start_in   (start_in_4_45),
       .swap_in   (swap_in_4_45),
       .op_in      (op_in_4_45),
       .pivot_in   (pivot_in_4_45),
       .start_out  (start_out_4_45),
       .swap_out   (swap_out_4_45),
       .data_out   (data_out_4_45),
       .op_out     (op_out_4_45),
       .pivot_out  (pivot_out_4_45),
       .r          (r_4_45)
     );

  // row 4, col 46

     reg start_in_4_46;
     wire start_out_4_46;

     reg swap_in_4_46;
     wire swap_out_4_46;

     reg [1:0] op_in_4_46;
     wire [1:0] op_out_4_46;

     wire r_4_46;

     reg data_in_4_46;
     wire data_out_4_46;

     reg pivot_in_4_46;
     wire pivot_out_4_46;

     always @(posedge clk) begin
         op_in_4_46 <= op_out_4_45;
         pivot_in_4_46 <= pivot_out_4_45;
         start_in_4_46 <= start_out_4_45;
         swap_in_4_46 <= swap_out_4_45;
     end

     always @(posedge clk) begin
         data_in_4_46 <= data_out_3_46;
     end
  
     processor_AB AB_4_46 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_46),
       .start_in   (start_in_4_46),
       .swap_in   (swap_in_4_46),
       .op_in      (op_in_4_46),
       .pivot_in   (pivot_in_4_46),
       .start_out  (start_out_4_46),
       .swap_out   (swap_out_4_46),
       .data_out   (data_out_4_46),
       .op_out     (op_out_4_46),
       .pivot_out  (pivot_out_4_46),
       .r          (r_4_46)
     );

  // row 4, col 47

     reg start_in_4_47;
     wire start_out_4_47;

     reg swap_in_4_47;
     wire swap_out_4_47;

     reg [1:0] op_in_4_47;
     wire [1:0] op_out_4_47;

     wire r_4_47;

     reg data_in_4_47;
     wire data_out_4_47;

     reg pivot_in_4_47;
     wire pivot_out_4_47;

     always @(posedge clk) begin
         op_in_4_47 <= op_out_4_46;
         pivot_in_4_47 <= pivot_out_4_46;
         start_in_4_47 <= start_out_4_46;
         swap_in_4_47 <= swap_out_4_46;
     end

     always @(posedge clk) begin
         data_in_4_47 <= data_out_3_47;
     end
  
     processor_AB AB_4_47 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_47),
       .start_in   (start_in_4_47),
       .swap_in   (swap_in_4_47),
       .op_in      (op_in_4_47),
       .pivot_in   (pivot_in_4_47),
       .start_out  (start_out_4_47),
       .swap_out   (swap_out_4_47),
       .data_out   (data_out_4_47),
       .op_out     (op_out_4_47),
       .pivot_out  (pivot_out_4_47),
       .r          (r_4_47)
     );

  // row 4, col 48

     reg start_in_4_48;
     wire start_out_4_48;

     reg swap_in_4_48;
     wire swap_out_4_48;

     reg [1:0] op_in_4_48;
     wire [1:0] op_out_4_48;

     wire r_4_48;

     reg data_in_4_48;
     wire data_out_4_48;

     reg pivot_in_4_48;
     wire pivot_out_4_48;

     always @(posedge clk) begin
         op_in_4_48 <= op_out_4_47;
         pivot_in_4_48 <= pivot_out_4_47;
         start_in_4_48 <= start_out_4_47;
         swap_in_4_48 <= swap_out_4_47;
     end

     always @(posedge clk) begin
         data_in_4_48 <= data_out_3_48;
     end
  
     processor_AB AB_4_48 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_48),
       .start_in   (start_in_4_48),
       .swap_in   (swap_in_4_48),
       .op_in      (op_in_4_48),
       .pivot_in   (pivot_in_4_48),
       .start_out  (start_out_4_48),
       .swap_out   (swap_out_4_48),
       .data_out   (data_out_4_48),
       .op_out     (op_out_4_48),
       .pivot_out  (pivot_out_4_48),
       .r          (r_4_48)
     );

  // row 4, col 49

     reg start_in_4_49;
     wire start_out_4_49;

     reg swap_in_4_49;
     wire swap_out_4_49;

     reg [1:0] op_in_4_49;
     wire [1:0] op_out_4_49;

     wire r_4_49;

     reg data_in_4_49;
     wire data_out_4_49;

     reg pivot_in_4_49;
     wire pivot_out_4_49;

     always @(posedge clk) begin
         op_in_4_49 <= op_out_4_48;
         pivot_in_4_49 <= pivot_out_4_48;
         start_in_4_49 <= start_out_4_48;
         swap_in_4_49 <= swap_out_4_48;
     end

     always @(posedge clk) begin
         data_in_4_49 <= data_out_3_49;
     end
  
     processor_AB AB_4_49 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_49),
       .start_in   (start_in_4_49),
       .swap_in   (swap_in_4_49),
       .op_in      (op_in_4_49),
       .pivot_in   (pivot_in_4_49),
       .start_out  (start_out_4_49),
       .swap_out   (swap_out_4_49),
       .data_out   (data_out_4_49),
       .op_out     (op_out_4_49),
       .pivot_out  (pivot_out_4_49),
       .r          (r_4_49)
     );

  // row 4, col 50

     reg start_in_4_50;
     wire start_out_4_50;

     reg swap_in_4_50;
     wire swap_out_4_50;

     reg [1:0] op_in_4_50;
     wire [1:0] op_out_4_50;

     wire r_4_50;

     reg data_in_4_50;
     wire data_out_4_50;

     reg pivot_in_4_50;
     wire pivot_out_4_50;

     always @(posedge clk) begin
         op_in_4_50 <= op_out_4_49;
         pivot_in_4_50 <= pivot_out_4_49;
         start_in_4_50 <= start_out_4_49;
         swap_in_4_50 <= swap_out_4_49;
     end

     always @(posedge clk) begin
         data_in_4_50 <= data_out_3_50;
     end
  
     processor_AB AB_4_50 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_50),
       .start_in   (start_in_4_50),
       .swap_in   (swap_in_4_50),
       .op_in      (op_in_4_50),
       .pivot_in   (pivot_in_4_50),
       .start_out  (start_out_4_50),
       .swap_out   (swap_out_4_50),
       .data_out   (data_out_4_50),
       .op_out     (op_out_4_50),
       .pivot_out  (pivot_out_4_50),
       .r          (r_4_50)
     );

  // row 4, col 51

     reg start_in_4_51;
     wire start_out_4_51;

     reg swap_in_4_51;
     wire swap_out_4_51;

     reg [1:0] op_in_4_51;
     wire [1:0] op_out_4_51;

     wire r_4_51;

     reg data_in_4_51;
     wire data_out_4_51;

     reg pivot_in_4_51;
     wire pivot_out_4_51;

     always @(posedge clk) begin
         op_in_4_51 <= op_out_4_50;
         pivot_in_4_51 <= pivot_out_4_50;
         start_in_4_51 <= start_out_4_50;
         swap_in_4_51 <= swap_out_4_50;
     end

     always @(posedge clk) begin
         data_in_4_51 <= data_out_3_51;
     end
  
     processor_AB AB_4_51 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_51),
       .start_in   (start_in_4_51),
       .swap_in   (swap_in_4_51),
       .op_in      (op_in_4_51),
       .pivot_in   (pivot_in_4_51),
       .start_out  (start_out_4_51),
       .swap_out   (swap_out_4_51),
       .data_out   (data_out_4_51),
       .op_out     (op_out_4_51),
       .pivot_out  (pivot_out_4_51),
       .r          (r_4_51)
     );

  // row 4, col 52

     reg start_in_4_52;
     wire start_out_4_52;

     reg swap_in_4_52;
     wire swap_out_4_52;

     reg [1:0] op_in_4_52;
     wire [1:0] op_out_4_52;

     wire r_4_52;

     reg data_in_4_52;
     wire data_out_4_52;

     reg pivot_in_4_52;
     wire pivot_out_4_52;

     always @(posedge clk) begin
         op_in_4_52 <= op_out_4_51;
         pivot_in_4_52 <= pivot_out_4_51;
         start_in_4_52 <= start_out_4_51;
         swap_in_4_52 <= swap_out_4_51;
     end

     always @(posedge clk) begin
         data_in_4_52 <= data_out_3_52;
     end
  
     processor_AB AB_4_52 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_52),
       .start_in   (start_in_4_52),
       .swap_in   (swap_in_4_52),
       .op_in      (op_in_4_52),
       .pivot_in   (pivot_in_4_52),
       .start_out  (start_out_4_52),
       .swap_out   (swap_out_4_52),
       .data_out   (data_out_4_52),
       .op_out     (op_out_4_52),
       .pivot_out  (pivot_out_4_52),
       .r          (r_4_52)
     );

  // row 4, col 53

     reg start_in_4_53;
     wire start_out_4_53;

     reg swap_in_4_53;
     wire swap_out_4_53;

     reg [1:0] op_in_4_53;
     wire [1:0] op_out_4_53;

     wire r_4_53;

     reg data_in_4_53;
     wire data_out_4_53;

     reg pivot_in_4_53;
     wire pivot_out_4_53;

     always @(posedge clk) begin
         op_in_4_53 <= op_out_4_52;
         pivot_in_4_53 <= pivot_out_4_52;
         start_in_4_53 <= start_out_4_52;
         swap_in_4_53 <= swap_out_4_52;
     end

     always @(posedge clk) begin
         data_in_4_53 <= data_out_3_53;
     end
  
     processor_AB AB_4_53 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_53),
       .start_in   (start_in_4_53),
       .swap_in   (swap_in_4_53),
       .op_in      (op_in_4_53),
       .pivot_in   (pivot_in_4_53),
       .start_out  (start_out_4_53),
       .swap_out   (swap_out_4_53),
       .data_out   (data_out_4_53),
       .op_out     (op_out_4_53),
       .pivot_out  (pivot_out_4_53),
       .r          (r_4_53)
     );

  // row 4, col 54

     reg start_in_4_54;
     wire start_out_4_54;

     reg swap_in_4_54;
     wire swap_out_4_54;

     reg [1:0] op_in_4_54;
     wire [1:0] op_out_4_54;

     wire r_4_54;

     reg data_in_4_54;
     wire data_out_4_54;

     reg pivot_in_4_54;
     wire pivot_out_4_54;

     always @(posedge clk) begin
         op_in_4_54 <= op_out_4_53;
         pivot_in_4_54 <= pivot_out_4_53;
         start_in_4_54 <= start_out_4_53;
         swap_in_4_54 <= swap_out_4_53;
     end

     always @(posedge clk) begin
         data_in_4_54 <= data_out_3_54;
     end
  
     processor_AB AB_4_54 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_54),
       .start_in   (start_in_4_54),
       .swap_in   (swap_in_4_54),
       .op_in      (op_in_4_54),
       .pivot_in   (pivot_in_4_54),
       .start_out  (start_out_4_54),
       .swap_out   (swap_out_4_54),
       .data_out   (data_out_4_54),
       .op_out     (op_out_4_54),
       .pivot_out  (pivot_out_4_54),
       .r          (r_4_54)
     );

  // row 4, col 55

     reg start_in_4_55;
     wire start_out_4_55;

     reg swap_in_4_55;
     wire swap_out_4_55;

     reg [1:0] op_in_4_55;
     wire [1:0] op_out_4_55;

     wire r_4_55;

     reg data_in_4_55;
     wire data_out_4_55;

     reg pivot_in_4_55;
     wire pivot_out_4_55;

     always @(posedge clk) begin
         op_in_4_55 <= op_out_4_54;
         pivot_in_4_55 <= pivot_out_4_54;
         start_in_4_55 <= start_out_4_54;
         swap_in_4_55 <= swap_out_4_54;
     end

     always @(posedge clk) begin
         data_in_4_55 <= data_out_3_55;
     end
  
     processor_AB AB_4_55 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_55),
       .start_in   (start_in_4_55),
       .swap_in   (swap_in_4_55),
       .op_in      (op_in_4_55),
       .pivot_in   (pivot_in_4_55),
       .start_out  (start_out_4_55),
       .swap_out   (swap_out_4_55),
       .data_out   (data_out_4_55),
       .op_out     (op_out_4_55),
       .pivot_out  (pivot_out_4_55),
       .r          (r_4_55)
     );

  // row 4, col 56

     reg start_in_4_56;
     wire start_out_4_56;

     reg swap_in_4_56;
     wire swap_out_4_56;

     reg [1:0] op_in_4_56;
     wire [1:0] op_out_4_56;

     wire r_4_56;

     reg data_in_4_56;
     wire data_out_4_56;

     reg pivot_in_4_56;
     wire pivot_out_4_56;

     always @(posedge clk) begin
         op_in_4_56 <= op_out_4_55;
         pivot_in_4_56 <= pivot_out_4_55;
         start_in_4_56 <= start_out_4_55;
         swap_in_4_56 <= swap_out_4_55;
     end

     always @(posedge clk) begin
         data_in_4_56 <= data_out_3_56;
     end
  
     processor_AB AB_4_56 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_56),
       .start_in   (start_in_4_56),
       .swap_in   (swap_in_4_56),
       .op_in      (op_in_4_56),
       .pivot_in   (pivot_in_4_56),
       .start_out  (start_out_4_56),
       .swap_out   (swap_out_4_56),
       .data_out   (data_out_4_56),
       .op_out     (op_out_4_56),
       .pivot_out  (pivot_out_4_56),
       .r          (r_4_56)
     );

  // row 4, col 57

     reg start_in_4_57;
     wire start_out_4_57;

     reg swap_in_4_57;
     wire swap_out_4_57;

     reg [1:0] op_in_4_57;
     wire [1:0] op_out_4_57;

     wire r_4_57;

     reg data_in_4_57;
     wire data_out_4_57;

     reg pivot_in_4_57;
     wire pivot_out_4_57;

     always @(posedge clk) begin
         op_in_4_57 <= op_out_4_56;
         pivot_in_4_57 <= pivot_out_4_56;
         start_in_4_57 <= start_out_4_56;
         swap_in_4_57 <= swap_out_4_56;
     end

     always @(posedge clk) begin
         data_in_4_57 <= data_out_3_57;
     end
  
     processor_AB AB_4_57 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_57),
       .start_in   (start_in_4_57),
       .swap_in   (swap_in_4_57),
       .op_in      (op_in_4_57),
       .pivot_in   (pivot_in_4_57),
       .start_out  (start_out_4_57),
       .swap_out   (swap_out_4_57),
       .data_out   (data_out_4_57),
       .op_out     (op_out_4_57),
       .pivot_out  (pivot_out_4_57),
       .r          (r_4_57)
     );

  // row 4, col 58

     reg start_in_4_58;
     wire start_out_4_58;

     reg swap_in_4_58;
     wire swap_out_4_58;

     reg [1:0] op_in_4_58;
     wire [1:0] op_out_4_58;

     wire r_4_58;

     reg data_in_4_58;
     wire data_out_4_58;

     reg pivot_in_4_58;
     wire pivot_out_4_58;

     always @(posedge clk) begin
         op_in_4_58 <= op_out_4_57;
         pivot_in_4_58 <= pivot_out_4_57;
         start_in_4_58 <= start_out_4_57;
         swap_in_4_58 <= swap_out_4_57;
     end

     always @(posedge clk) begin
         data_in_4_58 <= data_out_3_58;
     end
  
     processor_AB AB_4_58 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_58),
       .start_in   (start_in_4_58),
       .swap_in   (swap_in_4_58),
       .op_in      (op_in_4_58),
       .pivot_in   (pivot_in_4_58),
       .start_out  (start_out_4_58),
       .swap_out   (swap_out_4_58),
       .data_out   (data_out_4_58),
       .op_out     (op_out_4_58),
       .pivot_out  (pivot_out_4_58),
       .r          (r_4_58)
     );

  // row 4, col 59

     reg start_in_4_59;
     wire start_out_4_59;

     reg swap_in_4_59;
     wire swap_out_4_59;

     reg [1:0] op_in_4_59;
     wire [1:0] op_out_4_59;

     wire r_4_59;

     reg data_in_4_59;
     wire data_out_4_59;

     reg pivot_in_4_59;
     wire pivot_out_4_59;

     always @(posedge clk) begin
         op_in_4_59 <= op_out_4_58;
         pivot_in_4_59 <= pivot_out_4_58;
         start_in_4_59 <= start_out_4_58;
         swap_in_4_59 <= swap_out_4_58;
     end

     always @(posedge clk) begin
         data_in_4_59 <= data_out_3_59;
     end
  
     processor_AB AB_4_59 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_59),
       .start_in   (start_in_4_59),
       .swap_in   (swap_in_4_59),
       .op_in      (op_in_4_59),
       .pivot_in   (pivot_in_4_59),
       .start_out  (start_out_4_59),
       .swap_out   (swap_out_4_59),
       .data_out   (data_out_4_59),
       .op_out     (op_out_4_59),
       .pivot_out  (pivot_out_4_59),
       .r          (r_4_59)
     );

  // row 4, col 60

     reg start_in_4_60;
     wire start_out_4_60;

     reg swap_in_4_60;
     wire swap_out_4_60;

     reg [1:0] op_in_4_60;
     wire [1:0] op_out_4_60;

     wire r_4_60;

     reg data_in_4_60;
     wire data_out_4_60;

     reg pivot_in_4_60;
     wire pivot_out_4_60;

     always @(posedge clk) begin
         op_in_4_60 <= op_out_4_59;
         pivot_in_4_60 <= pivot_out_4_59;
         start_in_4_60 <= start_out_4_59;
         swap_in_4_60 <= swap_out_4_59;
     end

     always @(posedge clk) begin
         data_in_4_60 <= data_out_3_60;
     end
  
     processor_AB AB_4_60 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_60),
       .start_in   (start_in_4_60),
       .swap_in   (swap_in_4_60),
       .op_in      (op_in_4_60),
       .pivot_in   (pivot_in_4_60),
       .start_out  (start_out_4_60),
       .swap_out   (swap_out_4_60),
       .data_out   (data_out_4_60),
       .op_out     (op_out_4_60),
       .pivot_out  (pivot_out_4_60),
       .r          (r_4_60)
     );

  // row 4, col 61

     reg start_in_4_61;
     wire start_out_4_61;

     reg swap_in_4_61;
     wire swap_out_4_61;

     reg [1:0] op_in_4_61;
     wire [1:0] op_out_4_61;

     wire r_4_61;

     reg data_in_4_61;
     wire data_out_4_61;

     reg pivot_in_4_61;
     wire pivot_out_4_61;

     always @(posedge clk) begin
         op_in_4_61 <= op_out_4_60;
         pivot_in_4_61 <= pivot_out_4_60;
         start_in_4_61 <= start_out_4_60;
         swap_in_4_61 <= swap_out_4_60;
     end

     always @(posedge clk) begin
         data_in_4_61 <= data_out_3_61;
     end
  
     processor_AB AB_4_61 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_61),
       .start_in   (start_in_4_61),
       .swap_in   (swap_in_4_61),
       .op_in      (op_in_4_61),
       .pivot_in   (pivot_in_4_61),
       .start_out  (start_out_4_61),
       .swap_out   (swap_out_4_61),
       .data_out   (data_out_4_61),
       .op_out     (op_out_4_61),
       .pivot_out  (pivot_out_4_61),
       .r          (r_4_61)
     );

  // row 4, col 62

     reg start_in_4_62;
     wire start_out_4_62;

     reg swap_in_4_62;
     wire swap_out_4_62;

     reg [1:0] op_in_4_62;
     wire [1:0] op_out_4_62;

     wire r_4_62;

     reg data_in_4_62;
     wire data_out_4_62;

     reg pivot_in_4_62;
     wire pivot_out_4_62;

     always @(posedge clk) begin
         op_in_4_62 <= op_out_4_61;
         pivot_in_4_62 <= pivot_out_4_61;
         start_in_4_62 <= start_out_4_61;
         swap_in_4_62 <= swap_out_4_61;
     end

     always @(posedge clk) begin
         data_in_4_62 <= data_out_3_62;
     end
  
     processor_AB AB_4_62 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_62),
       .start_in   (start_in_4_62),
       .swap_in   (swap_in_4_62),
       .op_in      (op_in_4_62),
       .pivot_in   (pivot_in_4_62),
       .start_out  (start_out_4_62),
       .swap_out   (swap_out_4_62),
       .data_out   (data_out_4_62),
       .op_out     (op_out_4_62),
       .pivot_out  (pivot_out_4_62),
       .r          (r_4_62)
     );

  // row 4, col 63

     reg start_in_4_63;
     wire start_out_4_63;

     reg swap_in_4_63;
     wire swap_out_4_63;

     reg [1:0] op_in_4_63;
     wire [1:0] op_out_4_63;

     wire r_4_63;

     reg data_in_4_63;
     wire data_out_4_63;

     reg pivot_in_4_63;
     wire pivot_out_4_63;

     always @(posedge clk) begin
         op_in_4_63 <= op_out_4_62;
         pivot_in_4_63 <= pivot_out_4_62;
         start_in_4_63 <= start_out_4_62;
         swap_in_4_63 <= swap_out_4_62;
     end

     always @(posedge clk) begin
         data_in_4_63 <= data_out_3_63;
     end
  
     processor_AB AB_4_63 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_63),
       .start_in   (start_in_4_63),
       .swap_in   (swap_in_4_63),
       .op_in      (op_in_4_63),
       .pivot_in   (pivot_in_4_63),
       .start_out  (start_out_4_63),
       .swap_out   (swap_out_4_63),
       .data_out   (data_out_4_63),
       .op_out     (op_out_4_63),
       .pivot_out  (pivot_out_4_63),
       .r          (r_4_63)
     );

  // row 4, col 64

     reg start_in_4_64;
     wire start_out_4_64;

     reg swap_in_4_64;
     wire swap_out_4_64;

     reg [1:0] op_in_4_64;
     wire [1:0] op_out_4_64;

     wire r_4_64;

     reg data_in_4_64;
     wire data_out_4_64;

     reg pivot_in_4_64;
     wire pivot_out_4_64;

     always @(posedge clk) begin
         op_in_4_64 <= op_out_4_63;
         pivot_in_4_64 <= pivot_out_4_63;
         start_in_4_64 <= start_out_4_63;
         swap_in_4_64 <= swap_out_4_63;
     end

     always @(posedge clk) begin
         data_in_4_64 <= data_out_3_64;
     end
  
     processor_AB AB_4_64 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_64),
       .start_in   (start_in_4_64),
       .swap_in   (swap_in_4_64),
       .op_in      (op_in_4_64),
       .pivot_in   (pivot_in_4_64),
       .start_out  (start_out_4_64),
       .swap_out   (swap_out_4_64),
       .data_out   (data_out_4_64),
       .op_out     (op_out_4_64),
       .pivot_out  (pivot_out_4_64),
       .r          (r_4_64)
     );

  // row 4, col 65

     reg start_in_4_65;
     wire start_out_4_65;

     reg swap_in_4_65;
     wire swap_out_4_65;

     reg [1:0] op_in_4_65;
     wire [1:0] op_out_4_65;

     wire r_4_65;

     reg data_in_4_65;
     wire data_out_4_65;

     reg pivot_in_4_65;
     wire pivot_out_4_65;

     always @(posedge clk) begin
         op_in_4_65 <= op_out_4_64;
         pivot_in_4_65 <= pivot_out_4_64;
         start_in_4_65 <= start_out_4_64;
         swap_in_4_65 <= swap_out_4_64;
     end

     always @(posedge clk) begin
         data_in_4_65 <= data_out_3_65;
     end
  
     processor_AB AB_4_65 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_65),
       .start_in   (start_in_4_65),
       .swap_in   (swap_in_4_65),
       .op_in      (op_in_4_65),
       .pivot_in   (pivot_in_4_65),
       .start_out  (start_out_4_65),
       .swap_out   (swap_out_4_65),
       .data_out   (data_out_4_65),
       .op_out     (op_out_4_65),
       .pivot_out  (pivot_out_4_65),
       .r          (r_4_65)
     );

  // row 4, col 66

     reg start_in_4_66;
     wire start_out_4_66;

     reg swap_in_4_66;
     wire swap_out_4_66;

     reg [1:0] op_in_4_66;
     wire [1:0] op_out_4_66;

     wire r_4_66;

     reg data_in_4_66;
     wire data_out_4_66;

     reg pivot_in_4_66;
     wire pivot_out_4_66;

     always @(posedge clk) begin
         op_in_4_66 <= op_out_4_65;
         pivot_in_4_66 <= pivot_out_4_65;
         start_in_4_66 <= start_out_4_65;
         swap_in_4_66 <= swap_out_4_65;
     end

     always @(posedge clk) begin
         data_in_4_66 <= data_out_3_66;
     end
  
     processor_AB AB_4_66 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_66),
       .start_in   (start_in_4_66),
       .swap_in   (swap_in_4_66),
       .op_in      (op_in_4_66),
       .pivot_in   (pivot_in_4_66),
       .start_out  (start_out_4_66),
       .swap_out   (swap_out_4_66),
       .data_out   (data_out_4_66),
       .op_out     (op_out_4_66),
       .pivot_out  (pivot_out_4_66),
       .r          (r_4_66)
     );

  // row 4, col 67

     reg start_in_4_67;
     wire start_out_4_67;

     reg swap_in_4_67;
     wire swap_out_4_67;

     reg [1:0] op_in_4_67;
     wire [1:0] op_out_4_67;

     wire r_4_67;

     reg data_in_4_67;
     wire data_out_4_67;

     reg pivot_in_4_67;
     wire pivot_out_4_67;

     always @(posedge clk) begin
         op_in_4_67 <= op_out_4_66;
         pivot_in_4_67 <= pivot_out_4_66;
         start_in_4_67 <= start_out_4_66;
         swap_in_4_67 <= swap_out_4_66;
     end

     always @(posedge clk) begin
         data_in_4_67 <= data_out_3_67;
     end
  
     processor_AB AB_4_67 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_67),
       .start_in   (start_in_4_67),
       .swap_in   (swap_in_4_67),
       .op_in      (op_in_4_67),
       .pivot_in   (pivot_in_4_67),
       .start_out  (start_out_4_67),
       .swap_out   (swap_out_4_67),
       .data_out   (data_out_4_67),
       .op_out     (op_out_4_67),
       .pivot_out  (pivot_out_4_67),
       .r          (r_4_67)
     );

  // row 4, col 68

     reg start_in_4_68;
     wire start_out_4_68;

     reg swap_in_4_68;
     wire swap_out_4_68;

     reg [1:0] op_in_4_68;
     wire [1:0] op_out_4_68;

     wire r_4_68;

     reg data_in_4_68;
     wire data_out_4_68;

     reg pivot_in_4_68;
     wire pivot_out_4_68;

     always @(posedge clk) begin
         op_in_4_68 <= op_out_4_67;
         pivot_in_4_68 <= pivot_out_4_67;
         start_in_4_68 <= start_out_4_67;
         swap_in_4_68 <= swap_out_4_67;
     end

     always @(posedge clk) begin
         data_in_4_68 <= data_out_3_68;
     end
  
     processor_AB AB_4_68 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_68),
       .start_in   (start_in_4_68),
       .swap_in   (swap_in_4_68),
       .op_in      (op_in_4_68),
       .pivot_in   (pivot_in_4_68),
       .start_out  (start_out_4_68),
       .swap_out   (swap_out_4_68),
       .data_out   (data_out_4_68),
       .op_out     (op_out_4_68),
       .pivot_out  (pivot_out_4_68),
       .r          (r_4_68)
     );

  // row 4, col 69

     reg start_in_4_69;
     wire start_out_4_69;

     reg swap_in_4_69;
     wire swap_out_4_69;

     reg [1:0] op_in_4_69;
     wire [1:0] op_out_4_69;

     wire r_4_69;

     reg data_in_4_69;
     wire data_out_4_69;

     reg pivot_in_4_69;
     wire pivot_out_4_69;

     always @(posedge clk) begin
         op_in_4_69 <= op_out_4_68;
         pivot_in_4_69 <= pivot_out_4_68;
         start_in_4_69 <= start_out_4_68;
         swap_in_4_69 <= swap_out_4_68;
     end

     always @(posedge clk) begin
         data_in_4_69 <= data_out_3_69;
     end
  
     processor_AB AB_4_69 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_69),
       .start_in   (start_in_4_69),
       .swap_in   (swap_in_4_69),
       .op_in      (op_in_4_69),
       .pivot_in   (pivot_in_4_69),
       .start_out  (start_out_4_69),
       .swap_out   (swap_out_4_69),
       .data_out   (data_out_4_69),
       .op_out     (op_out_4_69),
       .pivot_out  (pivot_out_4_69),
       .r          (r_4_69)
     );

  // row 4, col 70

     reg start_in_4_70;
     wire start_out_4_70;

     reg swap_in_4_70;
     wire swap_out_4_70;

     reg [1:0] op_in_4_70;
     wire [1:0] op_out_4_70;

     wire r_4_70;

     reg data_in_4_70;
     wire data_out_4_70;

     reg pivot_in_4_70;
     wire pivot_out_4_70;

     always @(posedge clk) begin
         op_in_4_70 <= op_out_4_69;
         pivot_in_4_70 <= pivot_out_4_69;
         start_in_4_70 <= start_out_4_69;
         swap_in_4_70 <= swap_out_4_69;
     end

     always @(posedge clk) begin
         data_in_4_70 <= data_out_3_70;
     end
  
     processor_AB AB_4_70 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_70),
       .start_in   (start_in_4_70),
       .swap_in   (swap_in_4_70),
       .op_in      (op_in_4_70),
       .pivot_in   (pivot_in_4_70),
       .start_out  (start_out_4_70),
       .swap_out   (swap_out_4_70),
       .data_out   (data_out_4_70),
       .op_out     (op_out_4_70),
       .pivot_out  (pivot_out_4_70),
       .r          (r_4_70)
     );

  // row 4, col 71

     reg start_in_4_71;
     wire start_out_4_71;

     reg swap_in_4_71;
     wire swap_out_4_71;

     reg [1:0] op_in_4_71;
     wire [1:0] op_out_4_71;

     wire r_4_71;

     reg data_in_4_71;
     wire data_out_4_71;

     reg pivot_in_4_71;
     wire pivot_out_4_71;

     always @(posedge clk) begin
         op_in_4_71 <= op_out_4_70;
         pivot_in_4_71 <= pivot_out_4_70;
         start_in_4_71 <= start_out_4_70;
         swap_in_4_71 <= swap_out_4_70;
     end

     always @(posedge clk) begin
         data_in_4_71 <= data_out_3_71;
     end
  
     processor_AB AB_4_71 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_71),
       .start_in   (start_in_4_71),
       .swap_in   (swap_in_4_71),
       .op_in      (op_in_4_71),
       .pivot_in   (pivot_in_4_71),
       .start_out  (start_out_4_71),
       .swap_out   (swap_out_4_71),
       .data_out   (data_out_4_71),
       .op_out     (op_out_4_71),
       .pivot_out  (pivot_out_4_71),
       .r          (r_4_71)
     );

  // row 4, col 72

     reg start_in_4_72;
     wire start_out_4_72;

     reg swap_in_4_72;
     wire swap_out_4_72;

     reg [1:0] op_in_4_72;
     wire [1:0] op_out_4_72;

     wire r_4_72;

     reg data_in_4_72;
     wire data_out_4_72;

     reg pivot_in_4_72;
     wire pivot_out_4_72;

     always @(posedge clk) begin
         op_in_4_72 <= op_out_4_71;
         pivot_in_4_72 <= pivot_out_4_71;
         start_in_4_72 <= start_out_4_71;
         swap_in_4_72 <= swap_out_4_71;
     end

     always @(posedge clk) begin
         data_in_4_72 <= data_out_3_72;
     end
  
     processor_AB AB_4_72 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_72),
       .start_in   (start_in_4_72),
       .swap_in   (swap_in_4_72),
       .op_in      (op_in_4_72),
       .pivot_in   (pivot_in_4_72),
       .start_out  (start_out_4_72),
       .swap_out   (swap_out_4_72),
       .data_out   (data_out_4_72),
       .op_out     (op_out_4_72),
       .pivot_out  (pivot_out_4_72),
       .r          (r_4_72)
     );

  // row 4, col 73

     reg start_in_4_73;
     wire start_out_4_73;

     reg swap_in_4_73;
     wire swap_out_4_73;

     reg [1:0] op_in_4_73;
     wire [1:0] op_out_4_73;

     wire r_4_73;

     reg data_in_4_73;
     wire data_out_4_73;

     reg pivot_in_4_73;
     wire pivot_out_4_73;

     always @(posedge clk) begin
         op_in_4_73 <= op_out_4_72;
         pivot_in_4_73 <= pivot_out_4_72;
         start_in_4_73 <= start_out_4_72;
         swap_in_4_73 <= swap_out_4_72;
     end

     always @(posedge clk) begin
         data_in_4_73 <= data_out_3_73;
     end
  
     processor_AB AB_4_73 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_73),
       .start_in   (start_in_4_73),
       .swap_in   (swap_in_4_73),
       .op_in      (op_in_4_73),
       .pivot_in   (pivot_in_4_73),
       .start_out  (start_out_4_73),
       .swap_out   (swap_out_4_73),
       .data_out   (data_out_4_73),
       .op_out     (op_out_4_73),
       .pivot_out  (pivot_out_4_73),
       .r          (r_4_73)
     );

  // row 4, col 74

     reg start_in_4_74;
     wire start_out_4_74;

     reg swap_in_4_74;
     wire swap_out_4_74;

     reg [1:0] op_in_4_74;
     wire [1:0] op_out_4_74;

     wire r_4_74;

     reg data_in_4_74;
     wire data_out_4_74;

     reg pivot_in_4_74;
     wire pivot_out_4_74;

     always @(posedge clk) begin
         op_in_4_74 <= op_out_4_73;
         pivot_in_4_74 <= pivot_out_4_73;
         start_in_4_74 <= start_out_4_73;
         swap_in_4_74 <= swap_out_4_73;
     end

     always @(posedge clk) begin
         data_in_4_74 <= data_out_3_74;
     end
  
     processor_AB AB_4_74 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_74),
       .start_in   (start_in_4_74),
       .swap_in   (swap_in_4_74),
       .op_in      (op_in_4_74),
       .pivot_in   (pivot_in_4_74),
       .start_out  (start_out_4_74),
       .swap_out   (swap_out_4_74),
       .data_out   (data_out_4_74),
       .op_out     (op_out_4_74),
       .pivot_out  (pivot_out_4_74),
       .r          (r_4_74)
     );

  // row 4, col 75

     reg start_in_4_75;
     wire start_out_4_75;

     reg swap_in_4_75;
     wire swap_out_4_75;

     reg [1:0] op_in_4_75;
     wire [1:0] op_out_4_75;

     wire r_4_75;

     reg data_in_4_75;
     wire data_out_4_75;

     reg pivot_in_4_75;
     wire pivot_out_4_75;

     always @(posedge clk) begin
         op_in_4_75 <= op_out_4_74;
         pivot_in_4_75 <= pivot_out_4_74;
         start_in_4_75 <= start_out_4_74;
         swap_in_4_75 <= swap_out_4_74;
     end

     always @(posedge clk) begin
         data_in_4_75 <= data_out_3_75;
     end
  
     processor_AB AB_4_75 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_75),
       .start_in   (start_in_4_75),
       .swap_in   (swap_in_4_75),
       .op_in      (op_in_4_75),
       .pivot_in   (pivot_in_4_75),
       .start_out  (start_out_4_75),
       .swap_out   (swap_out_4_75),
       .data_out   (data_out_4_75),
       .op_out     (op_out_4_75),
       .pivot_out  (pivot_out_4_75),
       .r          (r_4_75)
     );

  // row 4, col 76

     reg start_in_4_76;
     wire start_out_4_76;

     reg swap_in_4_76;
     wire swap_out_4_76;

     reg [1:0] op_in_4_76;
     wire [1:0] op_out_4_76;

     wire r_4_76;

     reg data_in_4_76;
     wire data_out_4_76;

     reg pivot_in_4_76;
     wire pivot_out_4_76;

     always @(posedge clk) begin
         op_in_4_76 <= op_out_4_75;
         pivot_in_4_76 <= pivot_out_4_75;
         start_in_4_76 <= start_out_4_75;
         swap_in_4_76 <= swap_out_4_75;
     end

     always @(posedge clk) begin
         data_in_4_76 <= data_out_3_76;
     end
  
     processor_AB AB_4_76 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_76),
       .start_in   (start_in_4_76),
       .swap_in   (swap_in_4_76),
       .op_in      (op_in_4_76),
       .pivot_in   (pivot_in_4_76),
       .start_out  (start_out_4_76),
       .swap_out   (swap_out_4_76),
       .data_out   (data_out_4_76),
       .op_out     (op_out_4_76),
       .pivot_out  (pivot_out_4_76),
       .r          (r_4_76)
     );

  // row 4, col 77

     reg start_in_4_77;
     wire start_out_4_77;

     reg swap_in_4_77;
     wire swap_out_4_77;

     reg [1:0] op_in_4_77;
     wire [1:0] op_out_4_77;

     wire r_4_77;

     reg data_in_4_77;
     wire data_out_4_77;

     reg pivot_in_4_77;
     wire pivot_out_4_77;

     always @(posedge clk) begin
         op_in_4_77 <= op_out_4_76;
         pivot_in_4_77 <= pivot_out_4_76;
         start_in_4_77 <= start_out_4_76;
         swap_in_4_77 <= swap_out_4_76;
     end

     always @(posedge clk) begin
         data_in_4_77 <= data_out_3_77;
     end
  
     processor_AB AB_4_77 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_77),
       .start_in   (start_in_4_77),
       .swap_in   (swap_in_4_77),
       .op_in      (op_in_4_77),
       .pivot_in   (pivot_in_4_77),
       .start_out  (start_out_4_77),
       .swap_out   (swap_out_4_77),
       .data_out   (data_out_4_77),
       .op_out     (op_out_4_77),
       .pivot_out  (pivot_out_4_77),
       .r          (r_4_77)
     );

  // row 4, col 78

     reg start_in_4_78;
     wire start_out_4_78;

     reg swap_in_4_78;
     wire swap_out_4_78;

     reg [1:0] op_in_4_78;
     wire [1:0] op_out_4_78;

     wire r_4_78;

     reg data_in_4_78;
     wire data_out_4_78;

     reg pivot_in_4_78;
     wire pivot_out_4_78;

     always @(posedge clk) begin
         op_in_4_78 <= op_out_4_77;
         pivot_in_4_78 <= pivot_out_4_77;
         start_in_4_78 <= start_out_4_77;
         swap_in_4_78 <= swap_out_4_77;
     end

     always @(posedge clk) begin
         data_in_4_78 <= data_out_3_78;
     end
  
     processor_AB AB_4_78 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_78),
       .start_in   (start_in_4_78),
       .swap_in   (swap_in_4_78),
       .op_in      (op_in_4_78),
       .pivot_in   (pivot_in_4_78),
       .start_out  (start_out_4_78),
       .swap_out   (swap_out_4_78),
       .data_out   (data_out_4_78),
       .op_out     (op_out_4_78),
       .pivot_out  (pivot_out_4_78),
       .r          (r_4_78)
     );

  // row 4, col 79

     reg start_in_4_79;
     wire start_out_4_79;

     reg swap_in_4_79;
     wire swap_out_4_79;

     reg [1:0] op_in_4_79;
     wire [1:0] op_out_4_79;

     wire r_4_79;

     reg data_in_4_79;
     wire data_out_4_79;

     reg pivot_in_4_79;
     wire pivot_out_4_79;

     always @(posedge clk) begin
         op_in_4_79 <= op_out_4_78;
         pivot_in_4_79 <= pivot_out_4_78;
         start_in_4_79 <= start_out_4_78;
         swap_in_4_79 <= swap_out_4_78;
     end

     always @(posedge clk) begin
         data_in_4_79 <= data_out_3_79;
     end
  
     processor_AB AB_4_79 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_79),
       .start_in   (start_in_4_79),
       .swap_in   (swap_in_4_79),
       .op_in      (op_in_4_79),
       .pivot_in   (pivot_in_4_79),
       .start_out  (start_out_4_79),
       .swap_out   (swap_out_4_79),
       .data_out   (data_out_4_79),
       .op_out     (op_out_4_79),
       .pivot_out  (pivot_out_4_79),
       .r          (r_4_79)
     );

  // row 4, col 80

     reg start_in_4_80;
     wire start_out_4_80;

     reg swap_in_4_80;
     wire swap_out_4_80;

     reg [1:0] op_in_4_80;
     wire [1:0] op_out_4_80;

     wire r_4_80;

     reg data_in_4_80;
     wire data_out_4_80;

     reg pivot_in_4_80;
     wire pivot_out_4_80;

     always @(posedge clk) begin
         op_in_4_80 <= op_out_4_79;
         pivot_in_4_80 <= pivot_out_4_79;
         start_in_4_80 <= start_out_4_79;
         swap_in_4_80 <= swap_out_4_79;
     end

     always @(posedge clk) begin
         data_in_4_80 <= data_out_3_80;
     end
  
     processor_AB AB_4_80 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_80),
       .start_in   (start_in_4_80),
       .swap_in   (swap_in_4_80),
       .op_in      (op_in_4_80),
       .pivot_in   (pivot_in_4_80),
       .start_out  (start_out_4_80),
       .swap_out   (swap_out_4_80),
       .data_out   (data_out_4_80),
       .op_out     (op_out_4_80),
       .pivot_out  (pivot_out_4_80),
       .r          (r_4_80)
     );

  // row 4, col 81

     reg start_in_4_81;
     wire start_out_4_81;

     reg swap_in_4_81;
     wire swap_out_4_81;

     reg [1:0] op_in_4_81;
     wire [1:0] op_out_4_81;

     wire r_4_81;

     reg data_in_4_81;
     wire data_out_4_81;

     reg pivot_in_4_81;
     wire pivot_out_4_81;

     always @(posedge clk) begin
         op_in_4_81 <= op_out_4_80;
         pivot_in_4_81 <= pivot_out_4_80;
         start_in_4_81 <= start_out_4_80;
         swap_in_4_81 <= swap_out_4_80;
     end

     always @(posedge clk) begin
         data_in_4_81 <= data_out_3_81;
     end
  
     processor_AB AB_4_81 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_81),
       .start_in   (start_in_4_81),
       .swap_in   (swap_in_4_81),
       .op_in      (op_in_4_81),
       .pivot_in   (pivot_in_4_81),
       .start_out  (start_out_4_81),
       .swap_out   (swap_out_4_81),
       .data_out   (data_out_4_81),
       .op_out     (op_out_4_81),
       .pivot_out  (pivot_out_4_81),
       .r          (r_4_81)
     );

  // row 4, col 82

     reg start_in_4_82;
     wire start_out_4_82;

     reg swap_in_4_82;
     wire swap_out_4_82;

     reg [1:0] op_in_4_82;
     wire [1:0] op_out_4_82;

     wire r_4_82;

     reg data_in_4_82;
     wire data_out_4_82;

     reg pivot_in_4_82;
     wire pivot_out_4_82;

     always @(posedge clk) begin
         op_in_4_82 <= op_out_4_81;
         pivot_in_4_82 <= pivot_out_4_81;
         start_in_4_82 <= start_out_4_81;
         swap_in_4_82 <= swap_out_4_81;
     end

     always @(posedge clk) begin
         data_in_4_82 <= data_out_3_82;
     end
  
     processor_AB AB_4_82 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_82),
       .start_in   (start_in_4_82),
       .swap_in   (swap_in_4_82),
       .op_in      (op_in_4_82),
       .pivot_in   (pivot_in_4_82),
       .start_out  (start_out_4_82),
       .swap_out   (swap_out_4_82),
       .data_out   (data_out_4_82),
       .op_out     (op_out_4_82),
       .pivot_out  (pivot_out_4_82),
       .r          (r_4_82)
     );

  // row 4, col 83

     reg start_in_4_83;
     wire start_out_4_83;

     reg swap_in_4_83;
     wire swap_out_4_83;

     reg [1:0] op_in_4_83;
     wire [1:0] op_out_4_83;

     wire r_4_83;

     reg data_in_4_83;
     wire data_out_4_83;

     reg pivot_in_4_83;
     wire pivot_out_4_83;

     always @(posedge clk) begin
         op_in_4_83 <= op_out_4_82;
         pivot_in_4_83 <= pivot_out_4_82;
         start_in_4_83 <= start_out_4_82;
         swap_in_4_83 <= swap_out_4_82;
     end

     always @(posedge clk) begin
         data_in_4_83 <= data_out_3_83;
     end
  
     processor_AB AB_4_83 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_83),
       .start_in   (start_in_4_83),
       .swap_in   (swap_in_4_83),
       .op_in      (op_in_4_83),
       .pivot_in   (pivot_in_4_83),
       .start_out  (start_out_4_83),
       .swap_out   (swap_out_4_83),
       .data_out   (data_out_4_83),
       .op_out     (op_out_4_83),
       .pivot_out  (pivot_out_4_83),
       .r          (r_4_83)
     );

  // row 4, col 84

     reg start_in_4_84;
     wire start_out_4_84;

     reg swap_in_4_84;
     wire swap_out_4_84;

     reg [1:0] op_in_4_84;
     wire [1:0] op_out_4_84;

     wire r_4_84;

     reg data_in_4_84;
     wire data_out_4_84;

     reg pivot_in_4_84;
     wire pivot_out_4_84;

     always @(posedge clk) begin
         op_in_4_84 <= op_out_4_83;
         pivot_in_4_84 <= pivot_out_4_83;
         start_in_4_84 <= start_out_4_83;
         swap_in_4_84 <= swap_out_4_83;
     end

     always @(posedge clk) begin
         data_in_4_84 <= data_out_3_84;
     end
  
     processor_AB AB_4_84 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_84),
       .start_in   (start_in_4_84),
       .swap_in   (swap_in_4_84),
       .op_in      (op_in_4_84),
       .pivot_in   (pivot_in_4_84),
       .start_out  (start_out_4_84),
       .swap_out   (swap_out_4_84),
       .data_out   (data_out_4_84),
       .op_out     (op_out_4_84),
       .pivot_out  (pivot_out_4_84),
       .r          (r_4_84)
     );

  // row 4, col 85

     reg start_in_4_85;
     wire start_out_4_85;

     reg swap_in_4_85;
     wire swap_out_4_85;

     reg [1:0] op_in_4_85;
     wire [1:0] op_out_4_85;

     wire r_4_85;

     reg data_in_4_85;
     wire data_out_4_85;

     reg pivot_in_4_85;
     wire pivot_out_4_85;

     always @(posedge clk) begin
         op_in_4_85 <= op_out_4_84;
         pivot_in_4_85 <= pivot_out_4_84;
         start_in_4_85 <= start_out_4_84;
         swap_in_4_85 <= swap_out_4_84;
     end

     always @(posedge clk) begin
         data_in_4_85 <= data_out_3_85;
     end
  
     processor_AB AB_4_85 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_85),
       .start_in   (start_in_4_85),
       .swap_in   (swap_in_4_85),
       .op_in      (op_in_4_85),
       .pivot_in   (pivot_in_4_85),
       .start_out  (start_out_4_85),
       .swap_out   (swap_out_4_85),
       .data_out   (data_out_4_85),
       .op_out     (op_out_4_85),
       .pivot_out  (pivot_out_4_85),
       .r          (r_4_85)
     );

  // row 4, col 86

     reg start_in_4_86;
     wire start_out_4_86;

     reg swap_in_4_86;
     wire swap_out_4_86;

     reg [1:0] op_in_4_86;
     wire [1:0] op_out_4_86;

     wire r_4_86;

     reg data_in_4_86;
     wire data_out_4_86;

     reg pivot_in_4_86;
     wire pivot_out_4_86;

     always @(posedge clk) begin
         op_in_4_86 <= op_out_4_85;
         pivot_in_4_86 <= pivot_out_4_85;
         start_in_4_86 <= start_out_4_85;
         swap_in_4_86 <= swap_out_4_85;
     end

     always @(posedge clk) begin
         data_in_4_86 <= data_out_3_86;
     end
  
     processor_AB AB_4_86 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_86),
       .start_in   (start_in_4_86),
       .swap_in   (swap_in_4_86),
       .op_in      (op_in_4_86),
       .pivot_in   (pivot_in_4_86),
       .start_out  (start_out_4_86),
       .swap_out   (swap_out_4_86),
       .data_out   (data_out_4_86),
       .op_out     (op_out_4_86),
       .pivot_out  (pivot_out_4_86),
       .r          (r_4_86)
     );

  // row 4, col 87

     reg start_in_4_87;
     wire start_out_4_87;

     reg swap_in_4_87;
     wire swap_out_4_87;

     reg [1:0] op_in_4_87;
     wire [1:0] op_out_4_87;

     wire r_4_87;

     reg data_in_4_87;
     wire data_out_4_87;

     reg pivot_in_4_87;
     wire pivot_out_4_87;

     always @(posedge clk) begin
         op_in_4_87 <= op_out_4_86;
         pivot_in_4_87 <= pivot_out_4_86;
         start_in_4_87 <= start_out_4_86;
         swap_in_4_87 <= swap_out_4_86;
     end

     always @(posedge clk) begin
         data_in_4_87 <= data_out_3_87;
     end
  
     processor_AB AB_4_87 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_87),
       .start_in   (start_in_4_87),
       .swap_in   (swap_in_4_87),
       .op_in      (op_in_4_87),
       .pivot_in   (pivot_in_4_87),
       .start_out  (start_out_4_87),
       .swap_out   (swap_out_4_87),
       .data_out   (data_out_4_87),
       .op_out     (op_out_4_87),
       .pivot_out  (pivot_out_4_87),
       .r          (r_4_87)
     );

  // row 4, col 88

     reg start_in_4_88;
     wire start_out_4_88;

     reg swap_in_4_88;
     wire swap_out_4_88;

     reg [1:0] op_in_4_88;
     wire [1:0] op_out_4_88;

     wire r_4_88;

     reg data_in_4_88;
     wire data_out_4_88;

     reg pivot_in_4_88;
     wire pivot_out_4_88;

     always @(posedge clk) begin
         op_in_4_88 <= op_out_4_87;
         pivot_in_4_88 <= pivot_out_4_87;
         start_in_4_88 <= start_out_4_87;
         swap_in_4_88 <= swap_out_4_87;
     end

     always @(posedge clk) begin
         data_in_4_88 <= data_out_3_88;
     end
  
     processor_AB AB_4_88 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_88),
       .start_in   (start_in_4_88),
       .swap_in   (swap_in_4_88),
       .op_in      (op_in_4_88),
       .pivot_in   (pivot_in_4_88),
       .start_out  (start_out_4_88),
       .swap_out   (swap_out_4_88),
       .data_out   (data_out_4_88),
       .op_out     (op_out_4_88),
       .pivot_out  (pivot_out_4_88),
       .r          (r_4_88)
     );

  // row 4, col 89

     reg start_in_4_89;
     wire start_out_4_89;

     reg swap_in_4_89;
     wire swap_out_4_89;

     reg [1:0] op_in_4_89;
     wire [1:0] op_out_4_89;

     wire r_4_89;

     reg data_in_4_89;
     wire data_out_4_89;

     reg pivot_in_4_89;
     wire pivot_out_4_89;

     always @(posedge clk) begin
         op_in_4_89 <= op_out_4_88;
         pivot_in_4_89 <= pivot_out_4_88;
         start_in_4_89 <= start_out_4_88;
         swap_in_4_89 <= swap_out_4_88;
     end

     always @(posedge clk) begin
         data_in_4_89 <= data_out_3_89;
     end
  
     processor_AB AB_4_89 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_89),
       .start_in   (start_in_4_89),
       .swap_in   (swap_in_4_89),
       .op_in      (op_in_4_89),
       .pivot_in   (pivot_in_4_89),
       .start_out  (start_out_4_89),
       .swap_out   (swap_out_4_89),
       .data_out   (data_out_4_89),
       .op_out     (op_out_4_89),
       .pivot_out  (pivot_out_4_89),
       .r          (r_4_89)
     );

  // row 4, col 90

     reg start_in_4_90;
     wire start_out_4_90;

     reg swap_in_4_90;
     wire swap_out_4_90;

     reg [1:0] op_in_4_90;
     wire [1:0] op_out_4_90;

     wire r_4_90;

     reg data_in_4_90;
     wire data_out_4_90;

     reg pivot_in_4_90;
     wire pivot_out_4_90;

     always @(posedge clk) begin
         op_in_4_90 <= op_out_4_89;
         pivot_in_4_90 <= pivot_out_4_89;
         start_in_4_90 <= start_out_4_89;
         swap_in_4_90 <= swap_out_4_89;
     end

     always @(posedge clk) begin
         data_in_4_90 <= data_out_3_90;
     end
  
     processor_AB AB_4_90 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_90),
       .start_in   (start_in_4_90),
       .swap_in   (swap_in_4_90),
       .op_in      (op_in_4_90),
       .pivot_in   (pivot_in_4_90),
       .start_out  (start_out_4_90),
       .swap_out   (swap_out_4_90),
       .data_out   (data_out_4_90),
       .op_out     (op_out_4_90),
       .pivot_out  (pivot_out_4_90),
       .r          (r_4_90)
     );

  // row 4, col 91

     reg start_in_4_91;
     wire start_out_4_91;

     reg swap_in_4_91;
     wire swap_out_4_91;

     reg [1:0] op_in_4_91;
     wire [1:0] op_out_4_91;

     wire r_4_91;

     reg data_in_4_91;
     wire data_out_4_91;

     reg pivot_in_4_91;
     wire pivot_out_4_91;

     always @(posedge clk) begin
         op_in_4_91 <= op_out_4_90;
         pivot_in_4_91 <= pivot_out_4_90;
         start_in_4_91 <= start_out_4_90;
         swap_in_4_91 <= swap_out_4_90;
     end

     always @(posedge clk) begin
         data_in_4_91 <= data_out_3_91;
     end
  
     processor_AB AB_4_91 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_91),
       .start_in   (start_in_4_91),
       .swap_in   (swap_in_4_91),
       .op_in      (op_in_4_91),
       .pivot_in   (pivot_in_4_91),
       .start_out  (start_out_4_91),
       .swap_out   (swap_out_4_91),
       .data_out   (data_out_4_91),
       .op_out     (op_out_4_91),
       .pivot_out  (pivot_out_4_91),
       .r          (r_4_91)
     );

  // row 4, col 92

     reg start_in_4_92;
     wire start_out_4_92;

     reg swap_in_4_92;
     wire swap_out_4_92;

     reg [1:0] op_in_4_92;
     wire [1:0] op_out_4_92;

     wire r_4_92;

     reg data_in_4_92;
     wire data_out_4_92;

     reg pivot_in_4_92;
     wire pivot_out_4_92;

     always @(posedge clk) begin
         op_in_4_92 <= op_out_4_91;
         pivot_in_4_92 <= pivot_out_4_91;
         start_in_4_92 <= start_out_4_91;
         swap_in_4_92 <= swap_out_4_91;
     end

     always @(posedge clk) begin
         data_in_4_92 <= data_out_3_92;
     end
  
     processor_AB AB_4_92 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_92),
       .start_in   (start_in_4_92),
       .swap_in   (swap_in_4_92),
       .op_in      (op_in_4_92),
       .pivot_in   (pivot_in_4_92),
       .start_out  (start_out_4_92),
       .swap_out   (swap_out_4_92),
       .data_out   (data_out_4_92),
       .op_out     (op_out_4_92),
       .pivot_out  (pivot_out_4_92),
       .r          (r_4_92)
     );

  // row 4, col 93

     reg start_in_4_93;
     wire start_out_4_93;

     reg swap_in_4_93;
     wire swap_out_4_93;

     reg [1:0] op_in_4_93;
     wire [1:0] op_out_4_93;

     wire r_4_93;

     reg data_in_4_93;
     wire data_out_4_93;

     reg pivot_in_4_93;
     wire pivot_out_4_93;

     always @(posedge clk) begin
         op_in_4_93 <= op_out_4_92;
         pivot_in_4_93 <= pivot_out_4_92;
         start_in_4_93 <= start_out_4_92;
         swap_in_4_93 <= swap_out_4_92;
     end

     always @(posedge clk) begin
         data_in_4_93 <= data_out_3_93;
     end
  
     processor_AB AB_4_93 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_93),
       .start_in   (start_in_4_93),
       .swap_in   (swap_in_4_93),
       .op_in      (op_in_4_93),
       .pivot_in   (pivot_in_4_93),
       .start_out  (start_out_4_93),
       .swap_out   (swap_out_4_93),
       .data_out   (data_out_4_93),
       .op_out     (op_out_4_93),
       .pivot_out  (pivot_out_4_93),
       .r          (r_4_93)
     );

  // row 4, col 94

     reg start_in_4_94;
     wire start_out_4_94;

     reg swap_in_4_94;
     wire swap_out_4_94;

     reg [1:0] op_in_4_94;
     wire [1:0] op_out_4_94;

     wire r_4_94;

     reg data_in_4_94;
     wire data_out_4_94;

     reg pivot_in_4_94;
     wire pivot_out_4_94;

     always @(posedge clk) begin
         op_in_4_94 <= op_out_4_93;
         pivot_in_4_94 <= pivot_out_4_93;
         start_in_4_94 <= start_out_4_93;
         swap_in_4_94 <= swap_out_4_93;
     end

     always @(posedge clk) begin
         data_in_4_94 <= data_out_3_94;
     end
  
     processor_AB AB_4_94 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_94),
       .start_in   (start_in_4_94),
       .swap_in   (swap_in_4_94),
       .op_in      (op_in_4_94),
       .pivot_in   (pivot_in_4_94),
       .start_out  (start_out_4_94),
       .swap_out   (swap_out_4_94),
       .data_out   (data_out_4_94),
       .op_out     (op_out_4_94),
       .pivot_out  (pivot_out_4_94),
       .r          (r_4_94)
     );

  // row 4, col 95

     reg start_in_4_95;
     wire start_out_4_95;

     reg swap_in_4_95;
     wire swap_out_4_95;

     reg [1:0] op_in_4_95;
     wire [1:0] op_out_4_95;

     wire r_4_95;

     reg data_in_4_95;
     wire data_out_4_95;

     reg pivot_in_4_95;
     wire pivot_out_4_95;

     always @(posedge clk) begin
         op_in_4_95 <= op_out_4_94;
         pivot_in_4_95 <= pivot_out_4_94;
         start_in_4_95 <= start_out_4_94;
         swap_in_4_95 <= swap_out_4_94;
     end

     always @(posedge clk) begin
         data_in_4_95 <= data_out_3_95;
     end
  
     processor_AB AB_4_95 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_95),
       .start_in   (start_in_4_95),
       .swap_in   (swap_in_4_95),
       .op_in      (op_in_4_95),
       .pivot_in   (pivot_in_4_95),
       .start_out  (start_out_4_95),
       .swap_out   (swap_out_4_95),
       .data_out   (data_out_4_95),
       .op_out     (op_out_4_95),
       .pivot_out  (pivot_out_4_95),
       .r          (r_4_95)
     );

  // row 4, col 96

     reg start_in_4_96;
     wire start_out_4_96;

     reg swap_in_4_96;
     wire swap_out_4_96;

     reg [1:0] op_in_4_96;
     wire [1:0] op_out_4_96;

     wire r_4_96;

     reg data_in_4_96;
     wire data_out_4_96;

     reg pivot_in_4_96;
     wire pivot_out_4_96;

     always @(posedge clk) begin
         op_in_4_96 <= op_out_4_95;
         pivot_in_4_96 <= pivot_out_4_95;
         start_in_4_96 <= start_out_4_95;
         swap_in_4_96 <= swap_out_4_95;
     end

     always @(posedge clk) begin
         data_in_4_96 <= data_out_3_96;
     end
  
     processor_AB AB_4_96 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_96),
       .start_in   (start_in_4_96),
       .swap_in   (swap_in_4_96),
       .op_in      (op_in_4_96),
       .pivot_in   (pivot_in_4_96),
       .start_out  (start_out_4_96),
       .swap_out   (swap_out_4_96),
       .data_out   (data_out_4_96),
       .op_out     (op_out_4_96),
       .pivot_out  (pivot_out_4_96),
       .r          (r_4_96)
     );

  // row 4, col 97

     reg start_in_4_97;
     wire start_out_4_97;

     reg swap_in_4_97;
     wire swap_out_4_97;

     reg [1:0] op_in_4_97;
     wire [1:0] op_out_4_97;

     wire r_4_97;

     reg data_in_4_97;
     wire data_out_4_97;

     reg pivot_in_4_97;
     wire pivot_out_4_97;

     always @(posedge clk) begin
         op_in_4_97 <= op_out_4_96;
         pivot_in_4_97 <= pivot_out_4_96;
         start_in_4_97 <= start_out_4_96;
         swap_in_4_97 <= swap_out_4_96;
     end

     always @(posedge clk) begin
         data_in_4_97 <= data_out_3_97;
     end
  
     processor_AB AB_4_97 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_97),
       .start_in   (start_in_4_97),
       .swap_in   (swap_in_4_97),
       .op_in      (op_in_4_97),
       .pivot_in   (pivot_in_4_97),
       .start_out  (start_out_4_97),
       .swap_out   (swap_out_4_97),
       .data_out   (data_out_4_97),
       .op_out     (op_out_4_97),
       .pivot_out  (pivot_out_4_97),
       .r          (r_4_97)
     );

  // row 4, col 98

     reg start_in_4_98;
     wire start_out_4_98;

     reg swap_in_4_98;
     wire swap_out_4_98;

     reg [1:0] op_in_4_98;
     wire [1:0] op_out_4_98;

     wire r_4_98;

     reg data_in_4_98;
     wire data_out_4_98;

     reg pivot_in_4_98;
     wire pivot_out_4_98;

     always @(posedge clk) begin
         op_in_4_98 <= op_out_4_97;
         pivot_in_4_98 <= pivot_out_4_97;
         start_in_4_98 <= start_out_4_97;
         swap_in_4_98 <= swap_out_4_97;
     end

     always @(posedge clk) begin
         data_in_4_98 <= data_out_3_98;
     end
  
     processor_AB AB_4_98 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_98),
       .start_in   (start_in_4_98),
       .swap_in   (swap_in_4_98),
       .op_in      (op_in_4_98),
       .pivot_in   (pivot_in_4_98),
       .start_out  (start_out_4_98),
       .swap_out   (swap_out_4_98),
       .data_out   (data_out_4_98),
       .op_out     (op_out_4_98),
       .pivot_out  (pivot_out_4_98),
       .r          (r_4_98)
     );

  // row 4, col 99

     reg start_in_4_99;
     wire start_out_4_99;

     reg swap_in_4_99;
     wire swap_out_4_99;

     reg [1:0] op_in_4_99;
     wire [1:0] op_out_4_99;

     wire r_4_99;

     reg data_in_4_99;
     wire data_out_4_99;

     reg pivot_in_4_99;
     wire pivot_out_4_99;

     always @(posedge clk) begin
         op_in_4_99 <= op_out_4_98;
         pivot_in_4_99 <= pivot_out_4_98;
         start_in_4_99 <= start_out_4_98;
         swap_in_4_99 <= swap_out_4_98;
     end

     always @(posedge clk) begin
         data_in_4_99 <= data_out_3_99;
     end
  
     processor_AB AB_4_99 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_99),
       .start_in   (start_in_4_99),
       .swap_in   (swap_in_4_99),
       .op_in      (op_in_4_99),
       .pivot_in   (pivot_in_4_99),
       .start_out  (start_out_4_99),
       .swap_out   (swap_out_4_99),
       .data_out   (data_out_4_99),
       .op_out     (op_out_4_99),
       .pivot_out  (pivot_out_4_99),
       .r          (r_4_99)
     );

  // row 4, col 100

     reg start_in_4_100;
     wire start_out_4_100;

     reg swap_in_4_100;
     wire swap_out_4_100;

     reg [1:0] op_in_4_100;
     wire [1:0] op_out_4_100;

     wire r_4_100;

     reg data_in_4_100;
     wire data_out_4_100;

     reg pivot_in_4_100;
     wire pivot_out_4_100;

     always @(posedge clk) begin
         op_in_4_100 <= op_out_4_99;
         pivot_in_4_100 <= pivot_out_4_99;
         start_in_4_100 <= start_out_4_99;
         swap_in_4_100 <= swap_out_4_99;
     end

     always @(posedge clk) begin
         data_in_4_100 <= data_out_3_100;
     end
  
     processor_AB AB_4_100 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_100),
       .start_in   (start_in_4_100),
       .swap_in   (swap_in_4_100),
       .op_in      (op_in_4_100),
       .pivot_in   (pivot_in_4_100),
       .start_out  (start_out_4_100),
       .swap_out   (swap_out_4_100),
       .data_out   (data_out_4_100),
       .op_out     (op_out_4_100),
       .pivot_out  (pivot_out_4_100),
       .r          (r_4_100)
     );

  // row 4, col 101

     reg start_in_4_101;
     wire start_out_4_101;

     reg swap_in_4_101;
     wire swap_out_4_101;

     reg [1:0] op_in_4_101;
     wire [1:0] op_out_4_101;

     wire r_4_101;

     reg data_in_4_101;
     wire data_out_4_101;

     reg pivot_in_4_101;
     wire pivot_out_4_101;

     always @(posedge clk) begin
         op_in_4_101 <= op_out_4_100;
         pivot_in_4_101 <= pivot_out_4_100;
         start_in_4_101 <= start_out_4_100;
         swap_in_4_101 <= swap_out_4_100;
     end

     always @(posedge clk) begin
         data_in_4_101 <= data_out_3_101;
     end
  
     processor_AB AB_4_101 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_101),
       .start_in   (start_in_4_101),
       .swap_in   (swap_in_4_101),
       .op_in      (op_in_4_101),
       .pivot_in   (pivot_in_4_101),
       .start_out  (start_out_4_101),
       .swap_out   (swap_out_4_101),
       .data_out   (data_out_4_101),
       .op_out     (op_out_4_101),
       .pivot_out  (pivot_out_4_101),
       .r          (r_4_101)
     );

  // row 4, col 102

     reg start_in_4_102;
     wire start_out_4_102;

     reg swap_in_4_102;
     wire swap_out_4_102;

     reg [1:0] op_in_4_102;
     wire [1:0] op_out_4_102;

     wire r_4_102;

     reg data_in_4_102;
     wire data_out_4_102;

     reg pivot_in_4_102;
     wire pivot_out_4_102;

     always @(posedge clk) begin
         op_in_4_102 <= op_out_4_101;
         pivot_in_4_102 <= pivot_out_4_101;
         start_in_4_102 <= start_out_4_101;
         swap_in_4_102 <= swap_out_4_101;
     end

     always @(posedge clk) begin
         data_in_4_102 <= data_out_3_102;
     end
  
     processor_AB AB_4_102 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_102),
       .start_in   (start_in_4_102),
       .swap_in   (swap_in_4_102),
       .op_in      (op_in_4_102),
       .pivot_in   (pivot_in_4_102),
       .start_out  (start_out_4_102),
       .swap_out   (swap_out_4_102),
       .data_out   (data_out_4_102),
       .op_out     (op_out_4_102),
       .pivot_out  (pivot_out_4_102),
       .r          (r_4_102)
     );

  // row 4, col 103

     reg start_in_4_103;
     wire start_out_4_103;

     reg swap_in_4_103;
     wire swap_out_4_103;

     reg [1:0] op_in_4_103;
     wire [1:0] op_out_4_103;

     wire r_4_103;

     reg data_in_4_103;
     wire data_out_4_103;

     reg pivot_in_4_103;
     wire pivot_out_4_103;

     always @(posedge clk) begin
         op_in_4_103 <= op_out_4_102;
         pivot_in_4_103 <= pivot_out_4_102;
         start_in_4_103 <= start_out_4_102;
         swap_in_4_103 <= swap_out_4_102;
     end

     always @(posedge clk) begin
         data_in_4_103 <= data_out_3_103;
     end
  
     processor_AB AB_4_103 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_103),
       .start_in   (start_in_4_103),
       .swap_in   (swap_in_4_103),
       .op_in      (op_in_4_103),
       .pivot_in   (pivot_in_4_103),
       .start_out  (start_out_4_103),
       .swap_out   (swap_out_4_103),
       .data_out   (data_out_4_103),
       .op_out     (op_out_4_103),
       .pivot_out  (pivot_out_4_103),
       .r          (r_4_103)
     );

  // row 4, col 104

     reg start_in_4_104;
     wire start_out_4_104;

     reg swap_in_4_104;
     wire swap_out_4_104;

     reg [1:0] op_in_4_104;
     wire [1:0] op_out_4_104;

     wire r_4_104;

     reg data_in_4_104;
     wire data_out_4_104;

     reg pivot_in_4_104;
     wire pivot_out_4_104;

     always @(posedge clk) begin
         op_in_4_104 <= op_out_4_103;
         pivot_in_4_104 <= pivot_out_4_103;
         start_in_4_104 <= start_out_4_103;
         swap_in_4_104 <= swap_out_4_103;
     end

     always @(posedge clk) begin
         data_in_4_104 <= data_out_3_104;
     end
  
     processor_AB AB_4_104 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_104),
       .start_in   (start_in_4_104),
       .swap_in   (swap_in_4_104),
       .op_in      (op_in_4_104),
       .pivot_in   (pivot_in_4_104),
       .start_out  (start_out_4_104),
       .swap_out   (swap_out_4_104),
       .data_out   (data_out_4_104),
       .op_out     (op_out_4_104),
       .pivot_out  (pivot_out_4_104),
       .r          (r_4_104)
     );

  // row 4, col 105

     reg start_in_4_105;
     wire start_out_4_105;

     reg swap_in_4_105;
     wire swap_out_4_105;

     reg [1:0] op_in_4_105;
     wire [1:0] op_out_4_105;

     wire r_4_105;

     reg data_in_4_105;
     wire data_out_4_105;

     reg pivot_in_4_105;
     wire pivot_out_4_105;

     always @(posedge clk) begin
         op_in_4_105 <= op_out_4_104;
         pivot_in_4_105 <= pivot_out_4_104;
         start_in_4_105 <= start_out_4_104;
         swap_in_4_105 <= swap_out_4_104;
     end

     always @(posedge clk) begin
         data_in_4_105 <= data_out_3_105;
     end
  
     processor_AB AB_4_105 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_105),
       .start_in   (start_in_4_105),
       .swap_in   (swap_in_4_105),
       .op_in      (op_in_4_105),
       .pivot_in   (pivot_in_4_105),
       .start_out  (start_out_4_105),
       .swap_out   (swap_out_4_105),
       .data_out   (data_out_4_105),
       .op_out     (op_out_4_105),
       .pivot_out  (pivot_out_4_105),
       .r          (r_4_105)
     );

  // row 4, col 106

     reg start_in_4_106;
     wire start_out_4_106;

     reg swap_in_4_106;
     wire swap_out_4_106;

     reg [1:0] op_in_4_106;
     wire [1:0] op_out_4_106;

     wire r_4_106;

     reg data_in_4_106;
     wire data_out_4_106;

     reg pivot_in_4_106;
     wire pivot_out_4_106;

     always @(posedge clk) begin
         op_in_4_106 <= op_out_4_105;
         pivot_in_4_106 <= pivot_out_4_105;
         start_in_4_106 <= start_out_4_105;
         swap_in_4_106 <= swap_out_4_105;
     end

     always @(posedge clk) begin
         data_in_4_106 <= data_out_3_106;
     end
  
     processor_AB AB_4_106 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_106),
       .start_in   (start_in_4_106),
       .swap_in   (swap_in_4_106),
       .op_in      (op_in_4_106),
       .pivot_in   (pivot_in_4_106),
       .start_out  (start_out_4_106),
       .swap_out   (swap_out_4_106),
       .data_out   (data_out_4_106),
       .op_out     (op_out_4_106),
       .pivot_out  (pivot_out_4_106),
       .r          (r_4_106)
     );

  // row 4, col 107

     reg start_in_4_107;
     wire start_out_4_107;

     reg swap_in_4_107;
     wire swap_out_4_107;

     reg [1:0] op_in_4_107;
     wire [1:0] op_out_4_107;

     wire r_4_107;

     reg data_in_4_107;
     wire data_out_4_107;

     reg pivot_in_4_107;
     wire pivot_out_4_107;

     always @(posedge clk) begin
         op_in_4_107 <= op_out_4_106;
         pivot_in_4_107 <= pivot_out_4_106;
         start_in_4_107 <= start_out_4_106;
         swap_in_4_107 <= swap_out_4_106;
     end

     always @(posedge clk) begin
         data_in_4_107 <= data_out_3_107;
     end
  
     processor_AB AB_4_107 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_107),
       .start_in   (start_in_4_107),
       .swap_in   (swap_in_4_107),
       .op_in      (op_in_4_107),
       .pivot_in   (pivot_in_4_107),
       .start_out  (start_out_4_107),
       .swap_out   (swap_out_4_107),
       .data_out   (data_out_4_107),
       .op_out     (op_out_4_107),
       .pivot_out  (pivot_out_4_107),
       .r          (r_4_107)
     );

  // row 4, col 108

     reg start_in_4_108;
     wire start_out_4_108;

     reg swap_in_4_108;
     wire swap_out_4_108;

     reg [1:0] op_in_4_108;
     wire [1:0] op_out_4_108;

     wire r_4_108;

     reg data_in_4_108;
     wire data_out_4_108;

     reg pivot_in_4_108;
     wire pivot_out_4_108;

     always @(posedge clk) begin
         op_in_4_108 <= op_out_4_107;
         pivot_in_4_108 <= pivot_out_4_107;
         start_in_4_108 <= start_out_4_107;
         swap_in_4_108 <= swap_out_4_107;
     end

     always @(posedge clk) begin
         data_in_4_108 <= data_out_3_108;
     end
  
     processor_AB AB_4_108 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_108),
       .start_in   (start_in_4_108),
       .swap_in   (swap_in_4_108),
       .op_in      (op_in_4_108),
       .pivot_in   (pivot_in_4_108),
       .start_out  (start_out_4_108),
       .swap_out   (swap_out_4_108),
       .data_out   (data_out_4_108),
       .op_out     (op_out_4_108),
       .pivot_out  (pivot_out_4_108),
       .r          (r_4_108)
     );

  // row 4, col 109

     reg start_in_4_109;
     wire start_out_4_109;

     reg swap_in_4_109;
     wire swap_out_4_109;

     reg [1:0] op_in_4_109;
     wire [1:0] op_out_4_109;

     wire r_4_109;

     reg data_in_4_109;
     wire data_out_4_109;

     reg pivot_in_4_109;
     wire pivot_out_4_109;

     always @(posedge clk) begin
         op_in_4_109 <= op_out_4_108;
         pivot_in_4_109 <= pivot_out_4_108;
         start_in_4_109 <= start_out_4_108;
         swap_in_4_109 <= swap_out_4_108;
     end

     always @(posedge clk) begin
         data_in_4_109 <= data_out_3_109;
     end
  
     processor_AB AB_4_109 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_109),
       .start_in   (start_in_4_109),
       .swap_in   (swap_in_4_109),
       .op_in      (op_in_4_109),
       .pivot_in   (pivot_in_4_109),
       .start_out  (start_out_4_109),
       .swap_out   (swap_out_4_109),
       .data_out   (data_out_4_109),
       .op_out     (op_out_4_109),
       .pivot_out  (pivot_out_4_109),
       .r          (r_4_109)
     );

  // row 4, col 110

     reg start_in_4_110;
     wire start_out_4_110;

     reg swap_in_4_110;
     wire swap_out_4_110;

     reg [1:0] op_in_4_110;
     wire [1:0] op_out_4_110;

     wire r_4_110;

     reg data_in_4_110;
     wire data_out_4_110;

     reg pivot_in_4_110;
     wire pivot_out_4_110;

     always @(posedge clk) begin
         op_in_4_110 <= op_out_4_109;
         pivot_in_4_110 <= pivot_out_4_109;
         start_in_4_110 <= start_out_4_109;
         swap_in_4_110 <= swap_out_4_109;
     end

     always @(posedge clk) begin
         data_in_4_110 <= data_out_3_110;
     end
  
     processor_AB AB_4_110 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_110),
       .start_in   (start_in_4_110),
       .swap_in   (swap_in_4_110),
       .op_in      (op_in_4_110),
       .pivot_in   (pivot_in_4_110),
       .start_out  (start_out_4_110),
       .swap_out   (swap_out_4_110),
       .data_out   (data_out_4_110),
       .op_out     (op_out_4_110),
       .pivot_out  (pivot_out_4_110),
       .r          (r_4_110)
     );

  // row 4, col 111

     reg start_in_4_111;
     wire start_out_4_111;

     reg swap_in_4_111;
     wire swap_out_4_111;

     reg [1:0] op_in_4_111;
     wire [1:0] op_out_4_111;

     wire r_4_111;

     reg data_in_4_111;
     wire data_out_4_111;

     reg pivot_in_4_111;
     wire pivot_out_4_111;

     always @(posedge clk) begin
         op_in_4_111 <= op_out_4_110;
         pivot_in_4_111 <= pivot_out_4_110;
         start_in_4_111 <= start_out_4_110;
         swap_in_4_111 <= swap_out_4_110;
     end

     always @(posedge clk) begin
         data_in_4_111 <= data_out_3_111;
     end
  
     processor_AB AB_4_111 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_111),
       .start_in   (start_in_4_111),
       .swap_in   (swap_in_4_111),
       .op_in      (op_in_4_111),
       .pivot_in   (pivot_in_4_111),
       .start_out  (start_out_4_111),
       .swap_out   (swap_out_4_111),
       .data_out   (data_out_4_111),
       .op_out     (op_out_4_111),
       .pivot_out  (pivot_out_4_111),
       .r          (r_4_111)
     );

  // row 4, col 112

     reg start_in_4_112;
     wire start_out_4_112;

     reg swap_in_4_112;
     wire swap_out_4_112;

     reg [1:0] op_in_4_112;
     wire [1:0] op_out_4_112;

     wire r_4_112;

     reg data_in_4_112;
     wire data_out_4_112;

     reg pivot_in_4_112;
     wire pivot_out_4_112;

     always @(posedge clk) begin
         op_in_4_112 <= op_out_4_111;
         pivot_in_4_112 <= pivot_out_4_111;
         start_in_4_112 <= start_out_4_111;
         swap_in_4_112 <= swap_out_4_111;
     end

     always @(posedge clk) begin
         data_in_4_112 <= data_out_3_112;
     end
  
     processor_AB AB_4_112 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_112),
       .start_in   (start_in_4_112),
       .swap_in   (swap_in_4_112),
       .op_in      (op_in_4_112),
       .pivot_in   (pivot_in_4_112),
       .start_out  (start_out_4_112),
       .swap_out   (swap_out_4_112),
       .data_out   (data_out_4_112),
       .op_out     (op_out_4_112),
       .pivot_out  (pivot_out_4_112),
       .r          (r_4_112)
     );

  // row 4, col 113

     reg start_in_4_113;
     wire start_out_4_113;

     reg swap_in_4_113;
     wire swap_out_4_113;

     reg [1:0] op_in_4_113;
     wire [1:0] op_out_4_113;

     wire r_4_113;

     reg data_in_4_113;
     wire data_out_4_113;

     reg pivot_in_4_113;
     wire pivot_out_4_113;

     always @(posedge clk) begin
         op_in_4_113 <= op_out_4_112;
         pivot_in_4_113 <= pivot_out_4_112;
         start_in_4_113 <= start_out_4_112;
         swap_in_4_113 <= swap_out_4_112;
     end

     always @(posedge clk) begin
         data_in_4_113 <= data_out_3_113;
     end
  
     processor_AB AB_4_113 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_113),
       .start_in   (start_in_4_113),
       .swap_in   (swap_in_4_113),
       .op_in      (op_in_4_113),
       .pivot_in   (pivot_in_4_113),
       .start_out  (start_out_4_113),
       .swap_out   (swap_out_4_113),
       .data_out   (data_out_4_113),
       .op_out     (op_out_4_113),
       .pivot_out  (pivot_out_4_113),
       .r          (r_4_113)
     );

  // row 4, col 114

     reg start_in_4_114;
     wire start_out_4_114;

     reg swap_in_4_114;
     wire swap_out_4_114;

     reg [1:0] op_in_4_114;
     wire [1:0] op_out_4_114;

     wire r_4_114;

     reg data_in_4_114;
     wire data_out_4_114;

     reg pivot_in_4_114;
     wire pivot_out_4_114;

     always @(posedge clk) begin
         op_in_4_114 <= op_out_4_113;
         pivot_in_4_114 <= pivot_out_4_113;
         start_in_4_114 <= start_out_4_113;
         swap_in_4_114 <= swap_out_4_113;
     end

     always @(posedge clk) begin
         data_in_4_114 <= data_out_3_114;
     end
  
     processor_AB AB_4_114 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_114),
       .start_in   (start_in_4_114),
       .swap_in   (swap_in_4_114),
       .op_in      (op_in_4_114),
       .pivot_in   (pivot_in_4_114),
       .start_out  (start_out_4_114),
       .swap_out   (swap_out_4_114),
       .data_out   (data_out_4_114),
       .op_out     (op_out_4_114),
       .pivot_out  (pivot_out_4_114),
       .r          (r_4_114)
     );

  // row 4, col 115

     reg start_in_4_115;
     wire start_out_4_115;

     reg swap_in_4_115;
     wire swap_out_4_115;

     reg [1:0] op_in_4_115;
     wire [1:0] op_out_4_115;

     wire r_4_115;

     reg data_in_4_115;
     wire data_out_4_115;

     reg pivot_in_4_115;
     wire pivot_out_4_115;

     always @(posedge clk) begin
         op_in_4_115 <= op_out_4_114;
         pivot_in_4_115 <= pivot_out_4_114;
         start_in_4_115 <= start_out_4_114;
         swap_in_4_115 <= swap_out_4_114;
     end

     always @(posedge clk) begin
         data_in_4_115 <= data_out_3_115;
     end
  
     processor_AB AB_4_115 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_115),
       .start_in   (start_in_4_115),
       .swap_in   (swap_in_4_115),
       .op_in      (op_in_4_115),
       .pivot_in   (pivot_in_4_115),
       .start_out  (start_out_4_115),
       .swap_out   (swap_out_4_115),
       .data_out   (data_out_4_115),
       .op_out     (op_out_4_115),
       .pivot_out  (pivot_out_4_115),
       .r          (r_4_115)
     );

  // row 4, col 116

     reg start_in_4_116;
     wire start_out_4_116;

     reg swap_in_4_116;
     wire swap_out_4_116;

     reg [1:0] op_in_4_116;
     wire [1:0] op_out_4_116;

     wire r_4_116;

     reg data_in_4_116;
     wire data_out_4_116;

     reg pivot_in_4_116;
     wire pivot_out_4_116;

     always @(posedge clk) begin
         op_in_4_116 <= op_out_4_115;
         pivot_in_4_116 <= pivot_out_4_115;
         start_in_4_116 <= start_out_4_115;
         swap_in_4_116 <= swap_out_4_115;
     end

     always @(posedge clk) begin
         data_in_4_116 <= data_out_3_116;
     end
  
     processor_AB AB_4_116 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_116),
       .start_in   (start_in_4_116),
       .swap_in   (swap_in_4_116),
       .op_in      (op_in_4_116),
       .pivot_in   (pivot_in_4_116),
       .start_out  (start_out_4_116),
       .swap_out   (swap_out_4_116),
       .data_out   (data_out_4_116),
       .op_out     (op_out_4_116),
       .pivot_out  (pivot_out_4_116),
       .r          (r_4_116)
     );

  // row 4, col 117

     reg start_in_4_117;
     wire start_out_4_117;

     reg swap_in_4_117;
     wire swap_out_4_117;

     reg [1:0] op_in_4_117;
     wire [1:0] op_out_4_117;

     wire r_4_117;

     reg data_in_4_117;
     wire data_out_4_117;

     reg pivot_in_4_117;
     wire pivot_out_4_117;

     always @(posedge clk) begin
         op_in_4_117 <= op_out_4_116;
         pivot_in_4_117 <= pivot_out_4_116;
         start_in_4_117 <= start_out_4_116;
         swap_in_4_117 <= swap_out_4_116;
     end

     always @(posedge clk) begin
         data_in_4_117 <= data_out_3_117;
     end
  
     processor_AB AB_4_117 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_117),
       .start_in   (start_in_4_117),
       .swap_in   (swap_in_4_117),
       .op_in      (op_in_4_117),
       .pivot_in   (pivot_in_4_117),
       .start_out  (start_out_4_117),
       .swap_out   (swap_out_4_117),
       .data_out   (data_out_4_117),
       .op_out     (op_out_4_117),
       .pivot_out  (pivot_out_4_117),
       .r          (r_4_117)
     );

  // row 4, col 118

     reg start_in_4_118;
     wire start_out_4_118;

     reg swap_in_4_118;
     wire swap_out_4_118;

     reg [1:0] op_in_4_118;
     wire [1:0] op_out_4_118;

     wire r_4_118;

     reg data_in_4_118;
     wire data_out_4_118;

     reg pivot_in_4_118;
     wire pivot_out_4_118;

     always @(posedge clk) begin
         op_in_4_118 <= op_out_4_117;
         pivot_in_4_118 <= pivot_out_4_117;
         start_in_4_118 <= start_out_4_117;
         swap_in_4_118 <= swap_out_4_117;
     end

     always @(posedge clk) begin
         data_in_4_118 <= data_out_3_118;
     end
  
     processor_AB AB_4_118 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_118),
       .start_in   (start_in_4_118),
       .swap_in   (swap_in_4_118),
       .op_in      (op_in_4_118),
       .pivot_in   (pivot_in_4_118),
       .start_out  (start_out_4_118),
       .swap_out   (swap_out_4_118),
       .data_out   (data_out_4_118),
       .op_out     (op_out_4_118),
       .pivot_out  (pivot_out_4_118),
       .r          (r_4_118)
     );

  // row 4, col 119

     reg start_in_4_119;
     wire start_out_4_119;

     reg swap_in_4_119;
     wire swap_out_4_119;

     reg [1:0] op_in_4_119;
     wire [1:0] op_out_4_119;

     wire r_4_119;

     reg data_in_4_119;
     wire data_out_4_119;

     reg pivot_in_4_119;
     wire pivot_out_4_119;

     always @(posedge clk) begin
         op_in_4_119 <= op_out_4_118;
         pivot_in_4_119 <= pivot_out_4_118;
         start_in_4_119 <= start_out_4_118;
         swap_in_4_119 <= swap_out_4_118;
     end

     always @(posedge clk) begin
         data_in_4_119 <= data_out_3_119;
     end
  
     processor_AB AB_4_119 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_119),
       .start_in   (start_in_4_119),
       .swap_in   (swap_in_4_119),
       .op_in      (op_in_4_119),
       .pivot_in   (pivot_in_4_119),
       .start_out  (start_out_4_119),
       .swap_out   (swap_out_4_119),
       .data_out   (data_out_4_119),
       .op_out     (op_out_4_119),
       .pivot_out  (pivot_out_4_119),
       .r          (r_4_119)
     );

  // row 4, col 120

     reg start_in_4_120;
     wire start_out_4_120;

     reg swap_in_4_120;
     wire swap_out_4_120;

     reg [1:0] op_in_4_120;
     wire [1:0] op_out_4_120;

     wire r_4_120;

     reg data_in_4_120;
     wire data_out_4_120;

     reg pivot_in_4_120;
     wire pivot_out_4_120;

     always @(posedge clk) begin
         op_in_4_120 <= op_out_4_119;
         pivot_in_4_120 <= pivot_out_4_119;
         start_in_4_120 <= start_out_4_119;
         swap_in_4_120 <= swap_out_4_119;
     end

     always @(posedge clk) begin
         data_in_4_120 <= data_out_3_120;
     end
  
     processor_AB AB_4_120 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_120),
       .start_in   (start_in_4_120),
       .swap_in   (swap_in_4_120),
       .op_in      (op_in_4_120),
       .pivot_in   (pivot_in_4_120),
       .start_out  (start_out_4_120),
       .swap_out   (swap_out_4_120),
       .data_out   (data_out_4_120),
       .op_out     (op_out_4_120),
       .pivot_out  (pivot_out_4_120),
       .r          (r_4_120)
     );

  // row 4, col 121

     reg start_in_4_121;
     wire start_out_4_121;

     reg swap_in_4_121;
     wire swap_out_4_121;

     reg [1:0] op_in_4_121;
     wire [1:0] op_out_4_121;

     wire r_4_121;

     reg data_in_4_121;
     wire data_out_4_121;

     reg pivot_in_4_121;
     wire pivot_out_4_121;

     always @(posedge clk) begin
         op_in_4_121 <= op_out_4_120;
         pivot_in_4_121 <= pivot_out_4_120;
         start_in_4_121 <= start_out_4_120;
         swap_in_4_121 <= swap_out_4_120;
     end

     always @(posedge clk) begin
         data_in_4_121 <= data_out_3_121;
     end
  
     processor_AB AB_4_121 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_121),
       .start_in   (start_in_4_121),
       .swap_in   (swap_in_4_121),
       .op_in      (op_in_4_121),
       .pivot_in   (pivot_in_4_121),
       .start_out  (start_out_4_121),
       .swap_out   (swap_out_4_121),
       .data_out   (data_out_4_121),
       .op_out     (op_out_4_121),
       .pivot_out  (pivot_out_4_121),
       .r          (r_4_121)
     );

  // row 4, col 122

     reg start_in_4_122;
     wire start_out_4_122;

     reg swap_in_4_122;
     wire swap_out_4_122;

     reg [1:0] op_in_4_122;
     wire [1:0] op_out_4_122;

     wire r_4_122;

     reg data_in_4_122;
     wire data_out_4_122;

     reg pivot_in_4_122;
     wire pivot_out_4_122;

     always @(posedge clk) begin
         op_in_4_122 <= op_out_4_121;
         pivot_in_4_122 <= pivot_out_4_121;
         start_in_4_122 <= start_out_4_121;
         swap_in_4_122 <= swap_out_4_121;
     end

     always @(posedge clk) begin
         data_in_4_122 <= data_out_3_122;
     end
  
     processor_AB AB_4_122 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_122),
       .start_in   (start_in_4_122),
       .swap_in   (swap_in_4_122),
       .op_in      (op_in_4_122),
       .pivot_in   (pivot_in_4_122),
       .start_out  (start_out_4_122),
       .swap_out   (swap_out_4_122),
       .data_out   (data_out_4_122),
       .op_out     (op_out_4_122),
       .pivot_out  (pivot_out_4_122),
       .r          (r_4_122)
     );

  // row 4, col 123

     reg start_in_4_123;
     wire start_out_4_123;

     reg swap_in_4_123;
     wire swap_out_4_123;

     reg [1:0] op_in_4_123;
     wire [1:0] op_out_4_123;

     wire r_4_123;

     reg data_in_4_123;
     wire data_out_4_123;

     reg pivot_in_4_123;
     wire pivot_out_4_123;

     always @(posedge clk) begin
         op_in_4_123 <= op_out_4_122;
         pivot_in_4_123 <= pivot_out_4_122;
         start_in_4_123 <= start_out_4_122;
         swap_in_4_123 <= swap_out_4_122;
     end

     always @(posedge clk) begin
         data_in_4_123 <= data_out_3_123;
     end
  
     processor_AB AB_4_123 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_123),
       .start_in   (start_in_4_123),
       .swap_in   (swap_in_4_123),
       .op_in      (op_in_4_123),
       .pivot_in   (pivot_in_4_123),
       .start_out  (start_out_4_123),
       .swap_out   (swap_out_4_123),
       .data_out   (data_out_4_123),
       .op_out     (op_out_4_123),
       .pivot_out  (pivot_out_4_123),
       .r          (r_4_123)
     );

  // row 4, col 124

     reg start_in_4_124;
     wire start_out_4_124;

     reg swap_in_4_124;
     wire swap_out_4_124;

     reg [1:0] op_in_4_124;
     wire [1:0] op_out_4_124;

     wire r_4_124;

     reg data_in_4_124;
     wire data_out_4_124;

     reg pivot_in_4_124;
     wire pivot_out_4_124;

     always @(posedge clk) begin
         op_in_4_124 <= op_out_4_123;
         pivot_in_4_124 <= pivot_out_4_123;
         start_in_4_124 <= start_out_4_123;
         swap_in_4_124 <= swap_out_4_123;
     end

     always @(posedge clk) begin
         data_in_4_124 <= data_out_3_124;
     end
  
     processor_AB AB_4_124 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_124),
       .start_in   (start_in_4_124),
       .swap_in   (swap_in_4_124),
       .op_in      (op_in_4_124),
       .pivot_in   (pivot_in_4_124),
       .start_out  (start_out_4_124),
       .swap_out   (swap_out_4_124),
       .data_out   (data_out_4_124),
       .op_out     (op_out_4_124),
       .pivot_out  (pivot_out_4_124),
       .r          (r_4_124)
     );

  // row 4, col 125

     reg start_in_4_125;
     wire start_out_4_125;

     reg swap_in_4_125;
     wire swap_out_4_125;

     reg [1:0] op_in_4_125;
     wire [1:0] op_out_4_125;

     wire r_4_125;

     reg data_in_4_125;
     wire data_out_4_125;

     reg pivot_in_4_125;
     wire pivot_out_4_125;

     always @(posedge clk) begin
         op_in_4_125 <= op_out_4_124;
         pivot_in_4_125 <= pivot_out_4_124;
         start_in_4_125 <= start_out_4_124;
         swap_in_4_125 <= swap_out_4_124;
     end

     always @(posedge clk) begin
         data_in_4_125 <= data_out_3_125;
     end
  
     processor_AB AB_4_125 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_125),
       .start_in   (start_in_4_125),
       .swap_in   (swap_in_4_125),
       .op_in      (op_in_4_125),
       .pivot_in   (pivot_in_4_125),
       .start_out  (start_out_4_125),
       .swap_out   (swap_out_4_125),
       .data_out   (data_out_4_125),
       .op_out     (op_out_4_125),
       .pivot_out  (pivot_out_4_125),
       .r          (r_4_125)
     );

  // row 4, col 126

     reg start_in_4_126;
     wire start_out_4_126;

     reg swap_in_4_126;
     wire swap_out_4_126;

     reg [1:0] op_in_4_126;
     wire [1:0] op_out_4_126;

     wire r_4_126;

     reg data_in_4_126;
     wire data_out_4_126;

     reg pivot_in_4_126;
     wire pivot_out_4_126;

     always @(posedge clk) begin
         op_in_4_126 <= op_out_4_125;
         pivot_in_4_126 <= pivot_out_4_125;
         start_in_4_126 <= start_out_4_125;
         swap_in_4_126 <= swap_out_4_125;
     end

     always @(posedge clk) begin
         data_in_4_126 <= data_out_3_126;
     end
  
     processor_AB AB_4_126 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_126),
       .start_in   (start_in_4_126),
       .swap_in   (swap_in_4_126),
       .op_in      (op_in_4_126),
       .pivot_in   (pivot_in_4_126),
       .start_out  (start_out_4_126),
       .swap_out   (swap_out_4_126),
       .data_out   (data_out_4_126),
       .op_out     (op_out_4_126),
       .pivot_out  (pivot_out_4_126),
       .r          (r_4_126)
     );

  // row 4, col 127

     reg start_in_4_127;
     wire start_out_4_127;

     reg swap_in_4_127;
     wire swap_out_4_127;

     reg [1:0] op_in_4_127;
     wire [1:0] op_out_4_127;

     wire r_4_127;

     reg data_in_4_127;
     wire data_out_4_127;

     reg pivot_in_4_127;
     wire pivot_out_4_127;

     always @(posedge clk) begin
         op_in_4_127 <= op_out_4_126;
         pivot_in_4_127 <= pivot_out_4_126;
         start_in_4_127 <= start_out_4_126;
         swap_in_4_127 <= swap_out_4_126;
     end

     always @(posedge clk) begin
         data_in_4_127 <= data_out_3_127;
     end
  
     processor_AB AB_4_127 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_127),
       .start_in   (start_in_4_127),
       .swap_in   (swap_in_4_127),
       .op_in      (op_in_4_127),
       .pivot_in   (pivot_in_4_127),
       .start_out  (start_out_4_127),
       .swap_out   (swap_out_4_127),
       .data_out   (data_out_4_127),
       .op_out     (op_out_4_127),
       .pivot_out  (pivot_out_4_127),
       .r          (r_4_127)
     );

  // row 4, col 128

     reg start_in_4_128;
     wire start_out_4_128;

     reg swap_in_4_128;
     wire swap_out_4_128;

     reg [1:0] op_in_4_128;
     wire [1:0] op_out_4_128;

     wire r_4_128;

     reg data_in_4_128;
     wire data_out_4_128;

     reg pivot_in_4_128;
     wire pivot_out_4_128;

     always @(posedge clk) begin
         op_in_4_128 <= op_out_4_127;
         pivot_in_4_128 <= pivot_out_4_127;
         start_in_4_128 <= start_out_4_127;
         swap_in_4_128 <= swap_out_4_127;
     end

     always @(posedge clk) begin
         data_in_4_128 <= data_out_3_128;
     end
  
     processor_AB AB_4_128 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_128),
       .start_in   (start_in_4_128),
       .swap_in   (swap_in_4_128),
       .op_in      (op_in_4_128),
       .pivot_in   (pivot_in_4_128),
       .start_out  (start_out_4_128),
       .swap_out   (swap_out_4_128),
       .data_out   (data_out_4_128),
       .op_out     (op_out_4_128),
       .pivot_out  (pivot_out_4_128),
       .r          (r_4_128)
     );

  // row 4, col 129

     reg start_in_4_129;
     wire start_out_4_129;

     reg swap_in_4_129;
     wire swap_out_4_129;

     reg [1:0] op_in_4_129;
     wire [1:0] op_out_4_129;

     wire r_4_129;

     reg data_in_4_129;
     wire data_out_4_129;

     reg pivot_in_4_129;
     wire pivot_out_4_129;

     always @(posedge clk) begin
         op_in_4_129 <= op_out_4_128;
         pivot_in_4_129 <= pivot_out_4_128;
         start_in_4_129 <= start_out_4_128;
         swap_in_4_129 <= swap_out_4_128;
     end

     always @(posedge clk) begin
         data_in_4_129 <= data_out_3_129;
     end
  
     processor_AB AB_4_129 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_129),
       .start_in   (start_in_4_129),
       .swap_in   (swap_in_4_129),
       .op_in      (op_in_4_129),
       .pivot_in   (pivot_in_4_129),
       .start_out  (start_out_4_129),
       .swap_out   (swap_out_4_129),
       .data_out   (data_out_4_129),
       .op_out     (op_out_4_129),
       .pivot_out  (pivot_out_4_129),
       .r          (r_4_129)
     );

  // row 4, col 130

     reg start_in_4_130;
     wire start_out_4_130;

     reg swap_in_4_130;
     wire swap_out_4_130;

     reg [1:0] op_in_4_130;
     wire [1:0] op_out_4_130;

     wire r_4_130;

     reg data_in_4_130;
     wire data_out_4_130;

     reg pivot_in_4_130;
     wire pivot_out_4_130;

     always @(posedge clk) begin
         op_in_4_130 <= op_out_4_129;
         pivot_in_4_130 <= pivot_out_4_129;
         start_in_4_130 <= start_out_4_129;
         swap_in_4_130 <= swap_out_4_129;
     end

     always @(posedge clk) begin
         data_in_4_130 <= data_out_3_130;
     end
  
     processor_AB AB_4_130 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_130),
       .start_in   (start_in_4_130),
       .swap_in   (swap_in_4_130),
       .op_in      (op_in_4_130),
       .pivot_in   (pivot_in_4_130),
       .start_out  (start_out_4_130),
       .swap_out   (swap_out_4_130),
       .data_out   (data_out_4_130),
       .op_out     (op_out_4_130),
       .pivot_out  (pivot_out_4_130),
       .r          (r_4_130)
     );

  // row 4, col 131

     reg start_in_4_131;
     wire start_out_4_131;

     reg swap_in_4_131;
     wire swap_out_4_131;

     reg [1:0] op_in_4_131;
     wire [1:0] op_out_4_131;

     wire r_4_131;

     reg data_in_4_131;
     wire data_out_4_131;

     reg pivot_in_4_131;
     wire pivot_out_4_131;

     always @(posedge clk) begin
         op_in_4_131 <= op_out_4_130;
         pivot_in_4_131 <= pivot_out_4_130;
         start_in_4_131 <= start_out_4_130;
         swap_in_4_131 <= swap_out_4_130;
     end

     always @(posedge clk) begin
         data_in_4_131 <= data_out_3_131;
     end
  
     processor_AB AB_4_131 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_131),
       .start_in   (start_in_4_131),
       .swap_in   (swap_in_4_131),
       .op_in      (op_in_4_131),
       .pivot_in   (pivot_in_4_131),
       .start_out  (start_out_4_131),
       .swap_out   (swap_out_4_131),
       .data_out   (data_out_4_131),
       .op_out     (op_out_4_131),
       .pivot_out  (pivot_out_4_131),
       .r          (r_4_131)
     );

  // row 4, col 132

     reg start_in_4_132;
     wire start_out_4_132;

     reg swap_in_4_132;
     wire swap_out_4_132;

     reg [1:0] op_in_4_132;
     wire [1:0] op_out_4_132;

     wire r_4_132;

     reg data_in_4_132;
     wire data_out_4_132;

     reg pivot_in_4_132;
     wire pivot_out_4_132;

     always @(posedge clk) begin
         op_in_4_132 <= op_out_4_131;
         pivot_in_4_132 <= pivot_out_4_131;
         start_in_4_132 <= start_out_4_131;
         swap_in_4_132 <= swap_out_4_131;
     end

     always @(posedge clk) begin
         data_in_4_132 <= data_out_3_132;
     end
  
     processor_AB AB_4_132 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_132),
       .start_in   (start_in_4_132),
       .swap_in   (swap_in_4_132),
       .op_in      (op_in_4_132),
       .pivot_in   (pivot_in_4_132),
       .start_out  (start_out_4_132),
       .swap_out   (swap_out_4_132),
       .data_out   (data_out_4_132),
       .op_out     (op_out_4_132),
       .pivot_out  (pivot_out_4_132),
       .r          (r_4_132)
     );

  // row 4, col 133

     reg start_in_4_133;
     wire start_out_4_133;

     reg swap_in_4_133;
     wire swap_out_4_133;

     reg [1:0] op_in_4_133;
     wire [1:0] op_out_4_133;

     wire r_4_133;

     reg data_in_4_133;
     wire data_out_4_133;

     reg pivot_in_4_133;
     wire pivot_out_4_133;

     always @(posedge clk) begin
         op_in_4_133 <= op_out_4_132;
         pivot_in_4_133 <= pivot_out_4_132;
         start_in_4_133 <= start_out_4_132;
         swap_in_4_133 <= swap_out_4_132;
     end

     always @(posedge clk) begin
         data_in_4_133 <= data_out_3_133;
     end
  
     processor_AB AB_4_133 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_133),
       .start_in   (start_in_4_133),
       .swap_in   (swap_in_4_133),
       .op_in      (op_in_4_133),
       .pivot_in   (pivot_in_4_133),
       .start_out  (start_out_4_133),
       .swap_out   (swap_out_4_133),
       .data_out   (data_out_4_133),
       .op_out     (op_out_4_133),
       .pivot_out  (pivot_out_4_133),
       .r          (r_4_133)
     );

  // row 4, col 134

     reg start_in_4_134;
     wire start_out_4_134;

     reg swap_in_4_134;
     wire swap_out_4_134;

     reg [1:0] op_in_4_134;
     wire [1:0] op_out_4_134;

     wire r_4_134;

     reg data_in_4_134;
     wire data_out_4_134;

     reg pivot_in_4_134;
     wire pivot_out_4_134;

     always @(posedge clk) begin
         op_in_4_134 <= op_out_4_133;
         pivot_in_4_134 <= pivot_out_4_133;
         start_in_4_134 <= start_out_4_133;
         swap_in_4_134 <= swap_out_4_133;
     end

     always @(posedge clk) begin
         data_in_4_134 <= data_out_3_134;
     end
  
     processor_AB AB_4_134 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_134),
       .start_in   (start_in_4_134),
       .swap_in   (swap_in_4_134),
       .op_in      (op_in_4_134),
       .pivot_in   (pivot_in_4_134),
       .start_out  (start_out_4_134),
       .swap_out   (swap_out_4_134),
       .data_out   (data_out_4_134),
       .op_out     (op_out_4_134),
       .pivot_out  (pivot_out_4_134),
       .r          (r_4_134)
     );

  // row 4, col 135

     reg start_in_4_135;
     wire start_out_4_135;

     reg swap_in_4_135;
     wire swap_out_4_135;

     reg [1:0] op_in_4_135;
     wire [1:0] op_out_4_135;

     wire r_4_135;

     reg data_in_4_135;
     wire data_out_4_135;

     reg pivot_in_4_135;
     wire pivot_out_4_135;

     always @(posedge clk) begin
         op_in_4_135 <= op_out_4_134;
         pivot_in_4_135 <= pivot_out_4_134;
         start_in_4_135 <= start_out_4_134;
         swap_in_4_135 <= swap_out_4_134;
     end

     always @(posedge clk) begin
         data_in_4_135 <= data_out_3_135;
     end
  
     processor_AB AB_4_135 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_135),
       .start_in   (start_in_4_135),
       .swap_in   (swap_in_4_135),
       .op_in      (op_in_4_135),
       .pivot_in   (pivot_in_4_135),
       .start_out  (start_out_4_135),
       .swap_out   (swap_out_4_135),
       .data_out   (data_out_4_135),
       .op_out     (op_out_4_135),
       .pivot_out  (pivot_out_4_135),
       .r          (r_4_135)
     );

  // row 4, col 136

     reg start_in_4_136;
     wire start_out_4_136;

     reg swap_in_4_136;
     wire swap_out_4_136;

     reg [1:0] op_in_4_136;
     wire [1:0] op_out_4_136;

     wire r_4_136;

     reg data_in_4_136;
     wire data_out_4_136;

     reg pivot_in_4_136;
     wire pivot_out_4_136;

     always @(posedge clk) begin
         op_in_4_136 <= op_out_4_135;
         pivot_in_4_136 <= pivot_out_4_135;
         start_in_4_136 <= start_out_4_135;
         swap_in_4_136 <= swap_out_4_135;
     end

     always @(posedge clk) begin
         data_in_4_136 <= data_out_3_136;
     end
  
     processor_AB AB_4_136 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_136),
       .start_in   (start_in_4_136),
       .swap_in   (swap_in_4_136),
       .op_in      (op_in_4_136),
       .pivot_in   (pivot_in_4_136),
       .start_out  (start_out_4_136),
       .swap_out   (swap_out_4_136),
       .data_out   (data_out_4_136),
       .op_out     (op_out_4_136),
       .pivot_out  (pivot_out_4_136),
       .r          (r_4_136)
     );

  // row 4, col 137

     reg start_in_4_137;
     wire start_out_4_137;

     reg swap_in_4_137;
     wire swap_out_4_137;

     reg [1:0] op_in_4_137;
     wire [1:0] op_out_4_137;

     wire r_4_137;

     reg data_in_4_137;
     wire data_out_4_137;

     reg pivot_in_4_137;
     wire pivot_out_4_137;

     always @(posedge clk) begin
         op_in_4_137 <= op_out_4_136;
         pivot_in_4_137 <= pivot_out_4_136;
         start_in_4_137 <= start_out_4_136;
         swap_in_4_137 <= swap_out_4_136;
     end

     always @(posedge clk) begin
         data_in_4_137 <= data_out_3_137;
     end
  
     processor_AB AB_4_137 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_137),
       .start_in   (start_in_4_137),
       .swap_in   (swap_in_4_137),
       .op_in      (op_in_4_137),
       .pivot_in   (pivot_in_4_137),
       .start_out  (start_out_4_137),
       .swap_out   (swap_out_4_137),
       .data_out   (data_out_4_137),
       .op_out     (op_out_4_137),
       .pivot_out  (pivot_out_4_137),
       .r          (r_4_137)
     );

  // row 4, col 138

     reg start_in_4_138;
     wire start_out_4_138;

     reg swap_in_4_138;
     wire swap_out_4_138;

     reg [1:0] op_in_4_138;
     wire [1:0] op_out_4_138;

     wire r_4_138;

     reg data_in_4_138;
     wire data_out_4_138;

     reg pivot_in_4_138;
     wire pivot_out_4_138;

     always @(posedge clk) begin
         op_in_4_138 <= op_out_4_137;
         pivot_in_4_138 <= pivot_out_4_137;
         start_in_4_138 <= start_out_4_137;
         swap_in_4_138 <= swap_out_4_137;
     end

     always @(posedge clk) begin
         data_in_4_138 <= data_out_3_138;
     end
  
     processor_AB AB_4_138 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_138),
       .start_in   (start_in_4_138),
       .swap_in   (swap_in_4_138),
       .op_in      (op_in_4_138),
       .pivot_in   (pivot_in_4_138),
       .start_out  (start_out_4_138),
       .swap_out   (swap_out_4_138),
       .data_out   (data_out_4_138),
       .op_out     (op_out_4_138),
       .pivot_out  (pivot_out_4_138),
       .r          (r_4_138)
     );

  // row 4, col 139

     reg start_in_4_139;
     wire start_out_4_139;

     reg swap_in_4_139;
     wire swap_out_4_139;

     reg [1:0] op_in_4_139;
     wire [1:0] op_out_4_139;

     wire r_4_139;

     reg data_in_4_139;
     wire data_out_4_139;

     reg pivot_in_4_139;
     wire pivot_out_4_139;

     always @(posedge clk) begin
         op_in_4_139 <= op_out_4_138;
         pivot_in_4_139 <= pivot_out_4_138;
         start_in_4_139 <= start_out_4_138;
         swap_in_4_139 <= swap_out_4_138;
     end

     always @(posedge clk) begin
         data_in_4_139 <= data_out_3_139;
     end
  
     processor_AB AB_4_139 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_139),
       .start_in   (start_in_4_139),
       .swap_in   (swap_in_4_139),
       .op_in      (op_in_4_139),
       .pivot_in   (pivot_in_4_139),
       .start_out  (start_out_4_139),
       .swap_out   (swap_out_4_139),
       .data_out   (data_out_4_139),
       .op_out     (op_out_4_139),
       .pivot_out  (pivot_out_4_139),
       .r          (r_4_139)
     );

  // row 4, col 140

     reg start_in_4_140;
     wire start_out_4_140;

     reg swap_in_4_140;
     wire swap_out_4_140;

     reg [1:0] op_in_4_140;
     wire [1:0] op_out_4_140;

     wire r_4_140;

     reg data_in_4_140;
     wire data_out_4_140;

     reg pivot_in_4_140;
     wire pivot_out_4_140;

     always @(posedge clk) begin
         op_in_4_140 <= op_out_4_139;
         pivot_in_4_140 <= pivot_out_4_139;
         start_in_4_140 <= start_out_4_139;
         swap_in_4_140 <= swap_out_4_139;
     end

     always @(posedge clk) begin
         data_in_4_140 <= data_out_3_140;
     end
  
     processor_AB AB_4_140 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_140),
       .start_in   (start_in_4_140),
       .swap_in   (swap_in_4_140),
       .op_in      (op_in_4_140),
       .pivot_in   (pivot_in_4_140),
       .start_out  (start_out_4_140),
       .swap_out   (swap_out_4_140),
       .data_out   (data_out_4_140),
       .op_out     (op_out_4_140),
       .pivot_out  (pivot_out_4_140),
       .r          (r_4_140)
     );

  // row 4, col 141

     reg start_in_4_141;
     wire start_out_4_141;

     reg swap_in_4_141;
     wire swap_out_4_141;

     reg [1:0] op_in_4_141;
     wire [1:0] op_out_4_141;

     wire r_4_141;

     reg data_in_4_141;
     wire data_out_4_141;

     reg pivot_in_4_141;
     wire pivot_out_4_141;

     always @(posedge clk) begin
         op_in_4_141 <= op_out_4_140;
         pivot_in_4_141 <= pivot_out_4_140;
         start_in_4_141 <= start_out_4_140;
         swap_in_4_141 <= swap_out_4_140;
     end

     always @(posedge clk) begin
         data_in_4_141 <= data_out_3_141;
     end
  
     processor_AB AB_4_141 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_141),
       .start_in   (start_in_4_141),
       .swap_in   (swap_in_4_141),
       .op_in      (op_in_4_141),
       .pivot_in   (pivot_in_4_141),
       .start_out  (start_out_4_141),
       .swap_out   (swap_out_4_141),
       .data_out   (data_out_4_141),
       .op_out     (op_out_4_141),
       .pivot_out  (pivot_out_4_141),
       .r          (r_4_141)
     );

  // row 4, col 142

     reg start_in_4_142;
     wire start_out_4_142;

     reg swap_in_4_142;
     wire swap_out_4_142;

     reg [1:0] op_in_4_142;
     wire [1:0] op_out_4_142;

     wire r_4_142;

     reg data_in_4_142;
     wire data_out_4_142;

     reg pivot_in_4_142;
     wire pivot_out_4_142;

     always @(posedge clk) begin
         op_in_4_142 <= op_out_4_141;
         pivot_in_4_142 <= pivot_out_4_141;
         start_in_4_142 <= start_out_4_141;
         swap_in_4_142 <= swap_out_4_141;
     end

     always @(posedge clk) begin
         data_in_4_142 <= data_out_3_142;
     end
  
     processor_AB AB_4_142 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_142),
       .start_in   (start_in_4_142),
       .swap_in   (swap_in_4_142),
       .op_in      (op_in_4_142),
       .pivot_in   (pivot_in_4_142),
       .start_out  (start_out_4_142),
       .swap_out   (swap_out_4_142),
       .data_out   (data_out_4_142),
       .op_out     (op_out_4_142),
       .pivot_out  (pivot_out_4_142),
       .r          (r_4_142)
     );

  // row 4, col 143

     reg start_in_4_143;
     wire start_out_4_143;

     reg swap_in_4_143;
     wire swap_out_4_143;

     reg [1:0] op_in_4_143;
     wire [1:0] op_out_4_143;

     wire r_4_143;

     reg data_in_4_143;
     wire data_out_4_143;

     reg pivot_in_4_143;
     wire pivot_out_4_143;

     always @(posedge clk) begin
         op_in_4_143 <= op_out_4_142;
         pivot_in_4_143 <= pivot_out_4_142;
         start_in_4_143 <= start_out_4_142;
         swap_in_4_143 <= swap_out_4_142;
     end

     always @(posedge clk) begin
         data_in_4_143 <= data_out_3_143;
     end
  
     processor_AB AB_4_143 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_143),
       .start_in   (start_in_4_143),
       .swap_in   (swap_in_4_143),
       .op_in      (op_in_4_143),
       .pivot_in   (pivot_in_4_143),
       .start_out  (start_out_4_143),
       .swap_out   (swap_out_4_143),
       .data_out   (data_out_4_143),
       .op_out     (op_out_4_143),
       .pivot_out  (pivot_out_4_143),
       .r          (r_4_143)
     );

  // row 4, col 144

     reg start_in_4_144;
     wire start_out_4_144;

     reg swap_in_4_144;
     wire swap_out_4_144;

     reg [1:0] op_in_4_144;
     wire [1:0] op_out_4_144;

     wire r_4_144;

     reg data_in_4_144;
     wire data_out_4_144;

     reg pivot_in_4_144;
     wire pivot_out_4_144;

     always @(posedge clk) begin
         op_in_4_144 <= op_out_4_143;
         pivot_in_4_144 <= pivot_out_4_143;
         start_in_4_144 <= start_out_4_143;
         swap_in_4_144 <= swap_out_4_143;
     end

     always @(posedge clk) begin
         data_in_4_144 <= data_out_3_144;
     end
  
     processor_AB AB_4_144 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_144),
       .start_in   (start_in_4_144),
       .swap_in   (swap_in_4_144),
       .op_in      (op_in_4_144),
       .pivot_in   (pivot_in_4_144),
       .start_out  (start_out_4_144),
       .swap_out   (swap_out_4_144),
       .data_out   (data_out_4_144),
       .op_out     (op_out_4_144),
       .pivot_out  (pivot_out_4_144),
       .r          (r_4_144)
     );

  // row 4, col 145

     reg start_in_4_145;
     wire start_out_4_145;

     reg swap_in_4_145;
     wire swap_out_4_145;

     reg [1:0] op_in_4_145;
     wire [1:0] op_out_4_145;

     wire r_4_145;

     reg data_in_4_145;
     wire data_out_4_145;

     reg pivot_in_4_145;
     wire pivot_out_4_145;

     always @(posedge clk) begin
         op_in_4_145 <= op_out_4_144;
         pivot_in_4_145 <= pivot_out_4_144;
         start_in_4_145 <= start_out_4_144;
         swap_in_4_145 <= swap_out_4_144;
     end

     always @(posedge clk) begin
         data_in_4_145 <= data_out_3_145;
     end
  
     processor_AB AB_4_145 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_145),
       .start_in   (start_in_4_145),
       .swap_in   (swap_in_4_145),
       .op_in      (op_in_4_145),
       .pivot_in   (pivot_in_4_145),
       .start_out  (start_out_4_145),
       .swap_out   (swap_out_4_145),
       .data_out   (data_out_4_145),
       .op_out     (op_out_4_145),
       .pivot_out  (pivot_out_4_145),
       .r          (r_4_145)
     );

  // row 4, col 146

     reg start_in_4_146;
     wire start_out_4_146;

     reg swap_in_4_146;
     wire swap_out_4_146;

     reg [1:0] op_in_4_146;
     wire [1:0] op_out_4_146;

     wire r_4_146;

     reg data_in_4_146;
     wire data_out_4_146;

     reg pivot_in_4_146;
     wire pivot_out_4_146;

     always @(posedge clk) begin
         op_in_4_146 <= op_out_4_145;
         pivot_in_4_146 <= pivot_out_4_145;
         start_in_4_146 <= start_out_4_145;
         swap_in_4_146 <= swap_out_4_145;
     end

     always @(posedge clk) begin
         data_in_4_146 <= data_out_3_146;
     end
  
     processor_AB AB_4_146 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_146),
       .start_in   (start_in_4_146),
       .swap_in   (swap_in_4_146),
       .op_in      (op_in_4_146),
       .pivot_in   (pivot_in_4_146),
       .start_out  (start_out_4_146),
       .swap_out   (swap_out_4_146),
       .data_out   (data_out_4_146),
       .op_out     (op_out_4_146),
       .pivot_out  (pivot_out_4_146),
       .r          (r_4_146)
     );

  // row 4, col 147

     reg start_in_4_147;
     wire start_out_4_147;

     reg swap_in_4_147;
     wire swap_out_4_147;

     reg [1:0] op_in_4_147;
     wire [1:0] op_out_4_147;

     wire r_4_147;

     reg data_in_4_147;
     wire data_out_4_147;

     reg pivot_in_4_147;
     wire pivot_out_4_147;

     always @(posedge clk) begin
         op_in_4_147 <= op_out_4_146;
         pivot_in_4_147 <= pivot_out_4_146;
         start_in_4_147 <= start_out_4_146;
         swap_in_4_147 <= swap_out_4_146;
     end

     always @(posedge clk) begin
         data_in_4_147 <= data_out_3_147;
     end
  
     processor_AB AB_4_147 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_147),
       .start_in   (start_in_4_147),
       .swap_in   (swap_in_4_147),
       .op_in      (op_in_4_147),
       .pivot_in   (pivot_in_4_147),
       .start_out  (start_out_4_147),
       .swap_out   (swap_out_4_147),
       .data_out   (data_out_4_147),
       .op_out     (op_out_4_147),
       .pivot_out  (pivot_out_4_147),
       .r          (r_4_147)
     );

  // row 4, col 148

     reg start_in_4_148;
     wire start_out_4_148;

     reg swap_in_4_148;
     wire swap_out_4_148;

     reg [1:0] op_in_4_148;
     wire [1:0] op_out_4_148;

     wire r_4_148;

     reg data_in_4_148;
     wire data_out_4_148;

     reg pivot_in_4_148;
     wire pivot_out_4_148;

     always @(posedge clk) begin
         op_in_4_148 <= op_out_4_147;
         pivot_in_4_148 <= pivot_out_4_147;
         start_in_4_148 <= start_out_4_147;
         swap_in_4_148 <= swap_out_4_147;
     end

     always @(posedge clk) begin
         data_in_4_148 <= data_out_3_148;
     end
  
     processor_AB AB_4_148 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_148),
       .start_in   (start_in_4_148),
       .swap_in   (swap_in_4_148),
       .op_in      (op_in_4_148),
       .pivot_in   (pivot_in_4_148),
       .start_out  (start_out_4_148),
       .swap_out   (swap_out_4_148),
       .data_out   (data_out_4_148),
       .op_out     (op_out_4_148),
       .pivot_out  (pivot_out_4_148),
       .r          (r_4_148)
     );

  // row 4, col 149

     reg start_in_4_149;
     wire start_out_4_149;

     reg swap_in_4_149;
     wire swap_out_4_149;

     reg [1:0] op_in_4_149;
     wire [1:0] op_out_4_149;

     wire r_4_149;

     reg data_in_4_149;
     wire data_out_4_149;

     reg pivot_in_4_149;
     wire pivot_out_4_149;

     always @(posedge clk) begin
         op_in_4_149 <= op_out_4_148;
         pivot_in_4_149 <= pivot_out_4_148;
         start_in_4_149 <= start_out_4_148;
         swap_in_4_149 <= swap_out_4_148;
     end

     always @(posedge clk) begin
         data_in_4_149 <= data_out_3_149;
     end
  
     processor_AB AB_4_149 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_149),
       .start_in   (start_in_4_149),
       .swap_in   (swap_in_4_149),
       .op_in      (op_in_4_149),
       .pivot_in   (pivot_in_4_149),
       .start_out  (start_out_4_149),
       .swap_out   (swap_out_4_149),
       .data_out   (data_out_4_149),
       .op_out     (op_out_4_149),
       .pivot_out  (pivot_out_4_149),
       .r          (r_4_149)
     );

  // row 4, col 150

     reg start_in_4_150;
     wire start_out_4_150;

     reg swap_in_4_150;
     wire swap_out_4_150;

     reg [1:0] op_in_4_150;
     wire [1:0] op_out_4_150;

     wire r_4_150;

     reg data_in_4_150;
     wire data_out_4_150;

     reg pivot_in_4_150;
     wire pivot_out_4_150;

     always @(posedge clk) begin
         op_in_4_150 <= op_out_4_149;
         pivot_in_4_150 <= pivot_out_4_149;
         start_in_4_150 <= start_out_4_149;
         swap_in_4_150 <= swap_out_4_149;
     end

     always @(posedge clk) begin
         data_in_4_150 <= data_out_3_150;
     end
  
     processor_AB AB_4_150 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_150),
       .start_in   (start_in_4_150),
       .swap_in   (swap_in_4_150),
       .op_in      (op_in_4_150),
       .pivot_in   (pivot_in_4_150),
       .start_out  (start_out_4_150),
       .swap_out   (swap_out_4_150),
       .data_out   (data_out_4_150),
       .op_out     (op_out_4_150),
       .pivot_out  (pivot_out_4_150),
       .r          (r_4_150)
     );

  // row 4, col 151

     reg start_in_4_151;
     wire start_out_4_151;

     reg swap_in_4_151;
     wire swap_out_4_151;

     reg [1:0] op_in_4_151;
     wire [1:0] op_out_4_151;

     wire r_4_151;

     reg data_in_4_151;
     wire data_out_4_151;

     reg pivot_in_4_151;
     wire pivot_out_4_151;

     always @(posedge clk) begin
         op_in_4_151 <= op_out_4_150;
         pivot_in_4_151 <= pivot_out_4_150;
         start_in_4_151 <= start_out_4_150;
         swap_in_4_151 <= swap_out_4_150;
     end

     always @(posedge clk) begin
         data_in_4_151 <= data_out_3_151;
     end
  
     processor_AB AB_4_151 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_151),
       .start_in   (start_in_4_151),
       .swap_in   (swap_in_4_151),
       .op_in      (op_in_4_151),
       .pivot_in   (pivot_in_4_151),
       .start_out  (start_out_4_151),
       .swap_out   (swap_out_4_151),
       .data_out   (data_out_4_151),
       .op_out     (op_out_4_151),
       .pivot_out  (pivot_out_4_151),
       .r          (r_4_151)
     );

  // row 4, col 152

     reg start_in_4_152;
     wire start_out_4_152;

     reg swap_in_4_152;
     wire swap_out_4_152;

     reg [1:0] op_in_4_152;
     wire [1:0] op_out_4_152;

     wire r_4_152;

     reg data_in_4_152;
     wire data_out_4_152;

     reg pivot_in_4_152;
     wire pivot_out_4_152;

     always @(posedge clk) begin
         op_in_4_152 <= op_out_4_151;
         pivot_in_4_152 <= pivot_out_4_151;
         start_in_4_152 <= start_out_4_151;
         swap_in_4_152 <= swap_out_4_151;
     end

     always @(posedge clk) begin
         data_in_4_152 <= data_out_3_152;
     end
  
     processor_AB AB_4_152 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_152),
       .start_in   (start_in_4_152),
       .swap_in   (swap_in_4_152),
       .op_in      (op_in_4_152),
       .pivot_in   (pivot_in_4_152),
       .start_out  (start_out_4_152),
       .swap_out   (swap_out_4_152),
       .data_out   (data_out_4_152),
       .op_out     (op_out_4_152),
       .pivot_out  (pivot_out_4_152),
       .r          (r_4_152)
     );

  // row 4, col 153

     reg start_in_4_153;
     wire start_out_4_153;

     reg swap_in_4_153;
     wire swap_out_4_153;

     reg [1:0] op_in_4_153;
     wire [1:0] op_out_4_153;

     wire r_4_153;

     reg data_in_4_153;
     wire data_out_4_153;

     reg pivot_in_4_153;
     wire pivot_out_4_153;

     always @(posedge clk) begin
         op_in_4_153 <= op_out_4_152;
         pivot_in_4_153 <= pivot_out_4_152;
         start_in_4_153 <= start_out_4_152;
         swap_in_4_153 <= swap_out_4_152;
     end

     always @(posedge clk) begin
         data_in_4_153 <= data_out_3_153;
     end
  
     processor_AB AB_4_153 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_153),
       .start_in   (start_in_4_153),
       .swap_in   (swap_in_4_153),
       .op_in      (op_in_4_153),
       .pivot_in   (pivot_in_4_153),
       .start_out  (start_out_4_153),
       .swap_out   (swap_out_4_153),
       .data_out   (data_out_4_153),
       .op_out     (op_out_4_153),
       .pivot_out  (pivot_out_4_153),
       .r          (r_4_153)
     );

  // row 4, col 154

     reg start_in_4_154;
     wire start_out_4_154;

     reg swap_in_4_154;
     wire swap_out_4_154;

     reg [1:0] op_in_4_154;
     wire [1:0] op_out_4_154;

     wire r_4_154;

     reg data_in_4_154;
     wire data_out_4_154;

     reg pivot_in_4_154;
     wire pivot_out_4_154;

     always @(posedge clk) begin
         op_in_4_154 <= op_out_4_153;
         pivot_in_4_154 <= pivot_out_4_153;
         start_in_4_154 <= start_out_4_153;
         swap_in_4_154 <= swap_out_4_153;
     end

     always @(posedge clk) begin
         data_in_4_154 <= data_out_3_154;
     end
  
     processor_AB AB_4_154 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_154),
       .start_in   (start_in_4_154),
       .swap_in   (swap_in_4_154),
       .op_in      (op_in_4_154),
       .pivot_in   (pivot_in_4_154),
       .start_out  (start_out_4_154),
       .swap_out   (swap_out_4_154),
       .data_out   (data_out_4_154),
       .op_out     (op_out_4_154),
       .pivot_out  (pivot_out_4_154),
       .r          (r_4_154)
     );

  // row 4, col 155

     reg start_in_4_155;
     wire start_out_4_155;

     reg swap_in_4_155;
     wire swap_out_4_155;

     reg [1:0] op_in_4_155;
     wire [1:0] op_out_4_155;

     wire r_4_155;

     reg data_in_4_155;
     wire data_out_4_155;

     reg pivot_in_4_155;
     wire pivot_out_4_155;

     always @(posedge clk) begin
         op_in_4_155 <= op_out_4_154;
         pivot_in_4_155 <= pivot_out_4_154;
         start_in_4_155 <= start_out_4_154;
         swap_in_4_155 <= swap_out_4_154;
     end

     always @(posedge clk) begin
         data_in_4_155 <= data_out_3_155;
     end
  
     processor_AB AB_4_155 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_155),
       .start_in   (start_in_4_155),
       .swap_in   (swap_in_4_155),
       .op_in      (op_in_4_155),
       .pivot_in   (pivot_in_4_155),
       .start_out  (start_out_4_155),
       .swap_out   (swap_out_4_155),
       .data_out   (data_out_4_155),
       .op_out     (op_out_4_155),
       .pivot_out  (pivot_out_4_155),
       .r          (r_4_155)
     );

  // row 4, col 156

     reg start_in_4_156;
     wire start_out_4_156;

     reg swap_in_4_156;
     wire swap_out_4_156;

     reg [1:0] op_in_4_156;
     wire [1:0] op_out_4_156;

     wire r_4_156;

     reg data_in_4_156;
     wire data_out_4_156;

     reg pivot_in_4_156;
     wire pivot_out_4_156;

     always @(posedge clk) begin
         op_in_4_156 <= op_out_4_155;
         pivot_in_4_156 <= pivot_out_4_155;
         start_in_4_156 <= start_out_4_155;
         swap_in_4_156 <= swap_out_4_155;
     end

     always @(posedge clk) begin
         data_in_4_156 <= data_out_3_156;
     end
  
     processor_AB AB_4_156 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_156),
       .start_in   (start_in_4_156),
       .swap_in   (swap_in_4_156),
       .op_in      (op_in_4_156),
       .pivot_in   (pivot_in_4_156),
       .start_out  (start_out_4_156),
       .swap_out   (swap_out_4_156),
       .data_out   (data_out_4_156),
       .op_out     (op_out_4_156),
       .pivot_out  (pivot_out_4_156),
       .r          (r_4_156)
     );

  // row 4, col 157

     reg start_in_4_157;
     wire start_out_4_157;

     reg swap_in_4_157;
     wire swap_out_4_157;

     reg [1:0] op_in_4_157;
     wire [1:0] op_out_4_157;

     wire r_4_157;

     reg data_in_4_157;
     wire data_out_4_157;

     reg pivot_in_4_157;
     wire pivot_out_4_157;

     always @(posedge clk) begin
         op_in_4_157 <= op_out_4_156;
         pivot_in_4_157 <= pivot_out_4_156;
         start_in_4_157 <= start_out_4_156;
         swap_in_4_157 <= swap_out_4_156;
     end

     always @(posedge clk) begin
         data_in_4_157 <= data_out_3_157;
     end
  
     processor_AB AB_4_157 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_157),
       .start_in   (start_in_4_157),
       .swap_in   (swap_in_4_157),
       .op_in      (op_in_4_157),
       .pivot_in   (pivot_in_4_157),
       .start_out  (start_out_4_157),
       .swap_out   (swap_out_4_157),
       .data_out   (data_out_4_157),
       .op_out     (op_out_4_157),
       .pivot_out  (pivot_out_4_157),
       .r          (r_4_157)
     );

  // row 4, col 158

     reg start_in_4_158;
     wire start_out_4_158;

     reg swap_in_4_158;
     wire swap_out_4_158;

     reg [1:0] op_in_4_158;
     wire [1:0] op_out_4_158;

     wire r_4_158;

     reg data_in_4_158;
     wire data_out_4_158;

     reg pivot_in_4_158;
     wire pivot_out_4_158;

     always @(posedge clk) begin
         op_in_4_158 <= op_out_4_157;
         pivot_in_4_158 <= pivot_out_4_157;
         start_in_4_158 <= start_out_4_157;
         swap_in_4_158 <= swap_out_4_157;
     end

     always @(posedge clk) begin
         data_in_4_158 <= data_out_3_158;
     end
  
     processor_AB AB_4_158 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_158),
       .start_in   (start_in_4_158),
       .swap_in   (swap_in_4_158),
       .op_in      (op_in_4_158),
       .pivot_in   (pivot_in_4_158),
       .start_out  (start_out_4_158),
       .swap_out   (swap_out_4_158),
       .data_out   (data_out_4_158),
       .op_out     (op_out_4_158),
       .pivot_out  (pivot_out_4_158),
       .r          (r_4_158)
     );

  // row 4, col 159

     reg start_in_4_159;
     wire start_out_4_159;

     reg swap_in_4_159;
     wire swap_out_4_159;

     reg [1:0] op_in_4_159;
     wire [1:0] op_out_4_159;

     wire r_4_159;

     reg data_in_4_159;
     wire data_out_4_159;

     reg pivot_in_4_159;
     wire pivot_out_4_159;

     always @(posedge clk) begin
         op_in_4_159 <= op_out_4_158;
         pivot_in_4_159 <= pivot_out_4_158;
         start_in_4_159 <= start_out_4_158;
         swap_in_4_159 <= swap_out_4_158;
     end

     always @(posedge clk) begin
         data_in_4_159 <= data_out_3_159;
     end
  
     processor_AB AB_4_159 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_159),
       .start_in   (start_in_4_159),
       .swap_in   (swap_in_4_159),
       .op_in      (op_in_4_159),
       .pivot_in   (pivot_in_4_159),
       .start_out  (start_out_4_159),
       .swap_out   (swap_out_4_159),
       .data_out   (data_out_4_159),
       .op_out     (op_out_4_159),
       .pivot_out  (pivot_out_4_159),
       .r          (r_4_159)
     );

  // row 4, col 160

     reg start_in_4_160;
     wire start_out_4_160;

     reg swap_in_4_160;
     wire swap_out_4_160;

     reg [1:0] op_in_4_160;
     wire [1:0] op_out_4_160;

     wire r_4_160;

     reg data_in_4_160;
     wire data_out_4_160;

     reg pivot_in_4_160;
     wire pivot_out_4_160;

     always @(posedge clk) begin
         op_in_4_160 <= op_out_4_159;
         pivot_in_4_160 <= pivot_out_4_159;
         start_in_4_160 <= start_out_4_159;
         swap_in_4_160 <= swap_out_4_159;
     end

     always @(posedge clk) begin
         data_in_4_160 <= data_out_3_160;
     end
  
     processor_AB AB_4_160 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_160),
       .start_in   (start_in_4_160),
       .swap_in   (swap_in_4_160),
       .op_in      (op_in_4_160),
       .pivot_in   (pivot_in_4_160),
       .start_out  (start_out_4_160),
       .swap_out   (swap_out_4_160),
       .data_out   (data_out_4_160),
       .op_out     (op_out_4_160),
       .pivot_out  (pivot_out_4_160),
       .r          (r_4_160)
     );

  // row 4, col 161

     reg start_in_4_161;
     wire start_out_4_161;

     reg swap_in_4_161;
     wire swap_out_4_161;

     reg [1:0] op_in_4_161;
     wire [1:0] op_out_4_161;

     wire r_4_161;

     reg data_in_4_161;
     wire data_out_4_161;

     reg pivot_in_4_161;
     wire pivot_out_4_161;

     always @(posedge clk) begin
         op_in_4_161 <= op_out_4_160;
         pivot_in_4_161 <= pivot_out_4_160;
         start_in_4_161 <= start_out_4_160;
         swap_in_4_161 <= swap_out_4_160;
     end

     always @(posedge clk) begin
         data_in_4_161 <= data_out_3_161;
     end
  
     processor_AB AB_4_161 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_161),
       .start_in   (start_in_4_161),
       .swap_in   (swap_in_4_161),
       .op_in      (op_in_4_161),
       .pivot_in   (pivot_in_4_161),
       .start_out  (start_out_4_161),
       .swap_out   (swap_out_4_161),
       .data_out   (data_out_4_161),
       .op_out     (op_out_4_161),
       .pivot_out  (pivot_out_4_161),
       .r          (r_4_161)
     );

  // row 4, col 162

     reg start_in_4_162;
     wire start_out_4_162;

     reg swap_in_4_162;
     wire swap_out_4_162;

     reg [1:0] op_in_4_162;
     wire [1:0] op_out_4_162;

     wire r_4_162;

     reg data_in_4_162;
     wire data_out_4_162;

     reg pivot_in_4_162;
     wire pivot_out_4_162;

     always @(posedge clk) begin
         op_in_4_162 <= op_out_4_161;
         pivot_in_4_162 <= pivot_out_4_161;
         start_in_4_162 <= start_out_4_161;
         swap_in_4_162 <= swap_out_4_161;
     end

     always @(posedge clk) begin
         data_in_4_162 <= data_out_3_162;
     end
  
     processor_AB AB_4_162 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_162),
       .start_in   (start_in_4_162),
       .swap_in   (swap_in_4_162),
       .op_in      (op_in_4_162),
       .pivot_in   (pivot_in_4_162),
       .start_out  (start_out_4_162),
       .swap_out   (swap_out_4_162),
       .data_out   (data_out_4_162),
       .op_out     (op_out_4_162),
       .pivot_out  (pivot_out_4_162),
       .r          (r_4_162)
     );

  // row 4, col 163

     reg start_in_4_163;
     wire start_out_4_163;

     reg swap_in_4_163;
     wire swap_out_4_163;

     reg [1:0] op_in_4_163;
     wire [1:0] op_out_4_163;

     wire r_4_163;

     reg data_in_4_163;
     wire data_out_4_163;

     reg pivot_in_4_163;
     wire pivot_out_4_163;

     always @(posedge clk) begin
         op_in_4_163 <= op_out_4_162;
         pivot_in_4_163 <= pivot_out_4_162;
         start_in_4_163 <= start_out_4_162;
         swap_in_4_163 <= swap_out_4_162;
     end

     always @(posedge clk) begin
         data_in_4_163 <= data_out_3_163;
     end
  
     processor_AB AB_4_163 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_163),
       .start_in   (start_in_4_163),
       .swap_in   (swap_in_4_163),
       .op_in      (op_in_4_163),
       .pivot_in   (pivot_in_4_163),
       .start_out  (start_out_4_163),
       .swap_out   (swap_out_4_163),
       .data_out   (data_out_4_163),
       .op_out     (op_out_4_163),
       .pivot_out  (pivot_out_4_163),
       .r          (r_4_163)
     );

  // row 4, col 164

     reg start_in_4_164;
     wire start_out_4_164;

     reg swap_in_4_164;
     wire swap_out_4_164;

     reg [1:0] op_in_4_164;
     wire [1:0] op_out_4_164;

     wire r_4_164;

     reg data_in_4_164;
     wire data_out_4_164;

     reg pivot_in_4_164;
     wire pivot_out_4_164;

     always @(posedge clk) begin
         op_in_4_164 <= op_out_4_163;
         pivot_in_4_164 <= pivot_out_4_163;
         start_in_4_164 <= start_out_4_163;
         swap_in_4_164 <= swap_out_4_163;
     end

     always @(posedge clk) begin
         data_in_4_164 <= data_out_3_164;
     end
  
     processor_AB AB_4_164 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_164),
       .start_in   (start_in_4_164),
       .swap_in   (swap_in_4_164),
       .op_in      (op_in_4_164),
       .pivot_in   (pivot_in_4_164),
       .start_out  (start_out_4_164),
       .swap_out   (swap_out_4_164),
       .data_out   (data_out_4_164),
       .op_out     (op_out_4_164),
       .pivot_out  (pivot_out_4_164),
       .r          (r_4_164)
     );

  // row 4, col 165

     reg start_in_4_165;
     wire start_out_4_165;

     reg swap_in_4_165;
     wire swap_out_4_165;

     reg [1:0] op_in_4_165;
     wire [1:0] op_out_4_165;

     wire r_4_165;

     reg data_in_4_165;
     wire data_out_4_165;

     reg pivot_in_4_165;
     wire pivot_out_4_165;

     always @(posedge clk) begin
         op_in_4_165 <= op_out_4_164;
         pivot_in_4_165 <= pivot_out_4_164;
         start_in_4_165 <= start_out_4_164;
         swap_in_4_165 <= swap_out_4_164;
     end

     always @(posedge clk) begin
         data_in_4_165 <= data_out_3_165;
     end
  
     processor_AB AB_4_165 (
       .clk        (clk),
       .rst_b      (rst_b),
       .mode       (mode),
       .data_in    (data_in_4_165),
       .start_in   (start_in_4_165),
       .swap_in   (swap_in_4_165),
       .op_in      (op_in_4_165),
       .pivot_in   (pivot_in_4_165),
       .start_out  (start_out_4_165),
       .swap_out   (swap_out_4_165),
       .data_out   (data_out_4_165),
       .op_out     (op_out_4_165),
       .pivot_out  (pivot_out_4_165),
       .r          (r_4_165)
     );

  /////////////////////////////////////
  // outputs 

  wire [4:0] pivot_found;
  wire [165:0] row0, row1, row2, row3, row4;

  assign pivot_found = {r_0_0 | r_0_1 | r_0_2 | r_0_3 | r_0_4 | r_0_5 | r_0_6 | r_0_7 | r_0_8 | r_0_9 | r_0_10 | r_0_11 | r_0_12 | r_0_13 | r_0_14 | r_0_15 | r_0_16 | r_0_17 | r_0_18 | r_0_19 | r_0_20 | r_0_21 | r_0_22 | r_0_23 | r_0_24 | r_0_25 | r_0_26 | r_0_27 | r_0_28 | r_0_29 | r_0_30 | r_0_31 | r_0_32 | r_0_33 | r_0_34 | r_0_35 | r_0_36 | r_0_37 | r_0_38 | r_0_39 | r_0_40 | r_0_41 | r_0_42 | r_0_43 | r_0_44 | r_0_45 | r_0_46 | r_0_47 | r_0_48 | r_0_49 | r_0_50 | r_0_51 | r_0_52 | r_0_53 | r_0_54 | r_0_55 | r_0_56 | r_0_57 | r_0_58 | r_0_59 | r_0_60 | r_0_61 | r_0_62 | r_0_63 | r_0_64 | r_0_65 | r_0_66 | r_0_67 | r_0_68 | r_0_69 | r_0_70 | r_0_71 | r_0_72 | r_0_73 | r_0_74 | r_0_75 | r_0_76 | r_0_77 | r_0_78 | r_0_79 | r_0_80 | r_0_81 | r_0_82 | r_0_83 | r_0_84 | r_0_85 | r_0_86 | r_0_87 | r_0_88 | r_0_89 | r_0_90 | r_0_91 | r_0_92 | r_0_93 | r_0_94 | r_0_95 | r_0_96 | r_0_97 | r_0_98 | r_0_99 | r_0_100 | r_0_101 | r_0_102 | r_0_103 | r_0_104 | r_0_105 | r_0_106 | r_0_107 | r_0_108 | r_0_109 | r_0_110 | r_0_111 | r_0_112 | r_0_113 | r_0_114 | r_0_115 | r_0_116 | r_0_117 | r_0_118 | r_0_119 | r_0_120 | r_0_121 | r_0_122 | r_0_123 | r_0_124 | r_0_125 | r_0_126 | r_0_127 | r_0_128 | r_0_129 | r_0_130 | r_0_131 | r_0_132 | r_0_133 | r_0_134 | r_0_135 | r_0_136 | r_0_137 | r_0_138 | r_0_139 | r_0_140 | r_0_141 | r_0_142 | r_0_143 | r_0_144 | r_0_145 | r_0_146 | r_0_147 | r_0_148 | r_0_149 | r_0_150 | r_0_151 | r_0_152 | r_0_153 | r_0_154 | r_0_155 | r_0_156 | r_0_157 | r_0_158 | r_0_159 | r_0_160 | r_0_161 | r_0_162 | r_0_163 | r_0_164 | r_0_165, r_1_0 | r_1_1 | r_1_2 | r_1_3 | r_1_4 | r_1_5 | r_1_6 | r_1_7 | r_1_8 | r_1_9 | r_1_10 | r_1_11 | r_1_12 | r_1_13 | r_1_14 | r_1_15 | r_1_16 | r_1_17 | r_1_18 | r_1_19 | r_1_20 | r_1_21 | r_1_22 | r_1_23 | r_1_24 | r_1_25 | r_1_26 | r_1_27 | r_1_28 | r_1_29 | r_1_30 | r_1_31 | r_1_32 | r_1_33 | r_1_34 | r_1_35 | r_1_36 | r_1_37 | r_1_38 | r_1_39 | r_1_40 | r_1_41 | r_1_42 | r_1_43 | r_1_44 | r_1_45 | r_1_46 | r_1_47 | r_1_48 | r_1_49 | r_1_50 | r_1_51 | r_1_52 | r_1_53 | r_1_54 | r_1_55 | r_1_56 | r_1_57 | r_1_58 | r_1_59 | r_1_60 | r_1_61 | r_1_62 | r_1_63 | r_1_64 | r_1_65 | r_1_66 | r_1_67 | r_1_68 | r_1_69 | r_1_70 | r_1_71 | r_1_72 | r_1_73 | r_1_74 | r_1_75 | r_1_76 | r_1_77 | r_1_78 | r_1_79 | r_1_80 | r_1_81 | r_1_82 | r_1_83 | r_1_84 | r_1_85 | r_1_86 | r_1_87 | r_1_88 | r_1_89 | r_1_90 | r_1_91 | r_1_92 | r_1_93 | r_1_94 | r_1_95 | r_1_96 | r_1_97 | r_1_98 | r_1_99 | r_1_100 | r_1_101 | r_1_102 | r_1_103 | r_1_104 | r_1_105 | r_1_106 | r_1_107 | r_1_108 | r_1_109 | r_1_110 | r_1_111 | r_1_112 | r_1_113 | r_1_114 | r_1_115 | r_1_116 | r_1_117 | r_1_118 | r_1_119 | r_1_120 | r_1_121 | r_1_122 | r_1_123 | r_1_124 | r_1_125 | r_1_126 | r_1_127 | r_1_128 | r_1_129 | r_1_130 | r_1_131 | r_1_132 | r_1_133 | r_1_134 | r_1_135 | r_1_136 | r_1_137 | r_1_138 | r_1_139 | r_1_140 | r_1_141 | r_1_142 | r_1_143 | r_1_144 | r_1_145 | r_1_146 | r_1_147 | r_1_148 | r_1_149 | r_1_150 | r_1_151 | r_1_152 | r_1_153 | r_1_154 | r_1_155 | r_1_156 | r_1_157 | r_1_158 | r_1_159 | r_1_160 | r_1_161 | r_1_162 | r_1_163 | r_1_164 | r_1_165, r_2_0 | r_2_1 | r_2_2 | r_2_3 | r_2_4 | r_2_5 | r_2_6 | r_2_7 | r_2_8 | r_2_9 | r_2_10 | r_2_11 | r_2_12 | r_2_13 | r_2_14 | r_2_15 | r_2_16 | r_2_17 | r_2_18 | r_2_19 | r_2_20 | r_2_21 | r_2_22 | r_2_23 | r_2_24 | r_2_25 | r_2_26 | r_2_27 | r_2_28 | r_2_29 | r_2_30 | r_2_31 | r_2_32 | r_2_33 | r_2_34 | r_2_35 | r_2_36 | r_2_37 | r_2_38 | r_2_39 | r_2_40 | r_2_41 | r_2_42 | r_2_43 | r_2_44 | r_2_45 | r_2_46 | r_2_47 | r_2_48 | r_2_49 | r_2_50 | r_2_51 | r_2_52 | r_2_53 | r_2_54 | r_2_55 | r_2_56 | r_2_57 | r_2_58 | r_2_59 | r_2_60 | r_2_61 | r_2_62 | r_2_63 | r_2_64 | r_2_65 | r_2_66 | r_2_67 | r_2_68 | r_2_69 | r_2_70 | r_2_71 | r_2_72 | r_2_73 | r_2_74 | r_2_75 | r_2_76 | r_2_77 | r_2_78 | r_2_79 | r_2_80 | r_2_81 | r_2_82 | r_2_83 | r_2_84 | r_2_85 | r_2_86 | r_2_87 | r_2_88 | r_2_89 | r_2_90 | r_2_91 | r_2_92 | r_2_93 | r_2_94 | r_2_95 | r_2_96 | r_2_97 | r_2_98 | r_2_99 | r_2_100 | r_2_101 | r_2_102 | r_2_103 | r_2_104 | r_2_105 | r_2_106 | r_2_107 | r_2_108 | r_2_109 | r_2_110 | r_2_111 | r_2_112 | r_2_113 | r_2_114 | r_2_115 | r_2_116 | r_2_117 | r_2_118 | r_2_119 | r_2_120 | r_2_121 | r_2_122 | r_2_123 | r_2_124 | r_2_125 | r_2_126 | r_2_127 | r_2_128 | r_2_129 | r_2_130 | r_2_131 | r_2_132 | r_2_133 | r_2_134 | r_2_135 | r_2_136 | r_2_137 | r_2_138 | r_2_139 | r_2_140 | r_2_141 | r_2_142 | r_2_143 | r_2_144 | r_2_145 | r_2_146 | r_2_147 | r_2_148 | r_2_149 | r_2_150 | r_2_151 | r_2_152 | r_2_153 | r_2_154 | r_2_155 | r_2_156 | r_2_157 | r_2_158 | r_2_159 | r_2_160 | r_2_161 | r_2_162 | r_2_163 | r_2_164 | r_2_165, r_3_0 | r_3_1 | r_3_2 | r_3_3 | r_3_4 | r_3_5 | r_3_6 | r_3_7 | r_3_8 | r_3_9 | r_3_10 | r_3_11 | r_3_12 | r_3_13 | r_3_14 | r_3_15 | r_3_16 | r_3_17 | r_3_18 | r_3_19 | r_3_20 | r_3_21 | r_3_22 | r_3_23 | r_3_24 | r_3_25 | r_3_26 | r_3_27 | r_3_28 | r_3_29 | r_3_30 | r_3_31 | r_3_32 | r_3_33 | r_3_34 | r_3_35 | r_3_36 | r_3_37 | r_3_38 | r_3_39 | r_3_40 | r_3_41 | r_3_42 | r_3_43 | r_3_44 | r_3_45 | r_3_46 | r_3_47 | r_3_48 | r_3_49 | r_3_50 | r_3_51 | r_3_52 | r_3_53 | r_3_54 | r_3_55 | r_3_56 | r_3_57 | r_3_58 | r_3_59 | r_3_60 | r_3_61 | r_3_62 | r_3_63 | r_3_64 | r_3_65 | r_3_66 | r_3_67 | r_3_68 | r_3_69 | r_3_70 | r_3_71 | r_3_72 | r_3_73 | r_3_74 | r_3_75 | r_3_76 | r_3_77 | r_3_78 | r_3_79 | r_3_80 | r_3_81 | r_3_82 | r_3_83 | r_3_84 | r_3_85 | r_3_86 | r_3_87 | r_3_88 | r_3_89 | r_3_90 | r_3_91 | r_3_92 | r_3_93 | r_3_94 | r_3_95 | r_3_96 | r_3_97 | r_3_98 | r_3_99 | r_3_100 | r_3_101 | r_3_102 | r_3_103 | r_3_104 | r_3_105 | r_3_106 | r_3_107 | r_3_108 | r_3_109 | r_3_110 | r_3_111 | r_3_112 | r_3_113 | r_3_114 | r_3_115 | r_3_116 | r_3_117 | r_3_118 | r_3_119 | r_3_120 | r_3_121 | r_3_122 | r_3_123 | r_3_124 | r_3_125 | r_3_126 | r_3_127 | r_3_128 | r_3_129 | r_3_130 | r_3_131 | r_3_132 | r_3_133 | r_3_134 | r_3_135 | r_3_136 | r_3_137 | r_3_138 | r_3_139 | r_3_140 | r_3_141 | r_3_142 | r_3_143 | r_3_144 | r_3_145 | r_3_146 | r_3_147 | r_3_148 | r_3_149 | r_3_150 | r_3_151 | r_3_152 | r_3_153 | r_3_154 | r_3_155 | r_3_156 | r_3_157 | r_3_158 | r_3_159 | r_3_160 | r_3_161 | r_3_162 | r_3_163 | r_3_164 | r_3_165, r_4_0 | r_4_1 | r_4_2 | r_4_3 | r_4_4 | r_4_5 | r_4_6 | r_4_7 | r_4_8 | r_4_9 | r_4_10 | r_4_11 | r_4_12 | r_4_13 | r_4_14 | r_4_15 | r_4_16 | r_4_17 | r_4_18 | r_4_19 | r_4_20 | r_4_21 | r_4_22 | r_4_23 | r_4_24 | r_4_25 | r_4_26 | r_4_27 | r_4_28 | r_4_29 | r_4_30 | r_4_31 | r_4_32 | r_4_33 | r_4_34 | r_4_35 | r_4_36 | r_4_37 | r_4_38 | r_4_39 | r_4_40 | r_4_41 | r_4_42 | r_4_43 | r_4_44 | r_4_45 | r_4_46 | r_4_47 | r_4_48 | r_4_49 | r_4_50 | r_4_51 | r_4_52 | r_4_53 | r_4_54 | r_4_55 | r_4_56 | r_4_57 | r_4_58 | r_4_59 | r_4_60 | r_4_61 | r_4_62 | r_4_63 | r_4_64 | r_4_65 | r_4_66 | r_4_67 | r_4_68 | r_4_69 | r_4_70 | r_4_71 | r_4_72 | r_4_73 | r_4_74 | r_4_75 | r_4_76 | r_4_77 | r_4_78 | r_4_79 | r_4_80 | r_4_81 | r_4_82 | r_4_83 | r_4_84 | r_4_85 | r_4_86 | r_4_87 | r_4_88 | r_4_89 | r_4_90 | r_4_91 | r_4_92 | r_4_93 | r_4_94 | r_4_95 | r_4_96 | r_4_97 | r_4_98 | r_4_99 | r_4_100 | r_4_101 | r_4_102 | r_4_103 | r_4_104 | r_4_105 | r_4_106 | r_4_107 | r_4_108 | r_4_109 | r_4_110 | r_4_111 | r_4_112 | r_4_113 | r_4_114 | r_4_115 | r_4_116 | r_4_117 | r_4_118 | r_4_119 | r_4_120 | r_4_121 | r_4_122 | r_4_123 | r_4_124 | r_4_125 | r_4_126 | r_4_127 | r_4_128 | r_4_129 | r_4_130 | r_4_131 | r_4_132 | r_4_133 | r_4_134 | r_4_135 | r_4_136 | r_4_137 | r_4_138 | r_4_139 | r_4_140 | r_4_141 | r_4_142 | r_4_143 | r_4_144 | r_4_145 | r_4_146 | r_4_147 | r_4_148 | r_4_149 | r_4_150 | r_4_151 | r_4_152 | r_4_153 | r_4_154 | r_4_155 | r_4_156 | r_4_157 | r_4_158 | r_4_159 | r_4_160 | r_4_161 | r_4_162 | r_4_163 | r_4_164 | r_4_165};
  assign full_rank =  pivot_found == 5'b11111 ? 1'b1 : 1'b0;

  assign row0 = {r_0_0, r_0_1, r_0_2, r_0_3, r_0_4, r_0_5, r_0_6, r_0_7, r_0_8, r_0_9, r_0_10, r_0_11, r_0_12, r_0_13, r_0_14, r_0_15, r_0_16, r_0_17, r_0_18, r_0_19, r_0_20, r_0_21, r_0_22, r_0_23, r_0_24, r_0_25, r_0_26, r_0_27, r_0_28, r_0_29, r_0_30, r_0_31, r_0_32, r_0_33, r_0_34, r_0_35, r_0_36, r_0_37, r_0_38, r_0_39, r_0_40, r_0_41, r_0_42, r_0_43, r_0_44, r_0_45, r_0_46, r_0_47, r_0_48, r_0_49, r_0_50, r_0_51, r_0_52, r_0_53, r_0_54, r_0_55, r_0_56, r_0_57, r_0_58, r_0_59, r_0_60, r_0_61, r_0_62, r_0_63, r_0_64, r_0_65, r_0_66, r_0_67, r_0_68, r_0_69, r_0_70, r_0_71, r_0_72, r_0_73, r_0_74, r_0_75, r_0_76, r_0_77, r_0_78, r_0_79, r_0_80, r_0_81, r_0_82, r_0_83, r_0_84, r_0_85, r_0_86, r_0_87, r_0_88, r_0_89, r_0_90, r_0_91, r_0_92, r_0_93, r_0_94, r_0_95, r_0_96, r_0_97, r_0_98, r_0_99, r_0_100, r_0_101, r_0_102, r_0_103, r_0_104, r_0_105, r_0_106, r_0_107, r_0_108, r_0_109, r_0_110, r_0_111, r_0_112, r_0_113, r_0_114, r_0_115, r_0_116, r_0_117, r_0_118, r_0_119, r_0_120, r_0_121, r_0_122, r_0_123, r_0_124, r_0_125, r_0_126, r_0_127, r_0_128, r_0_129, r_0_130, r_0_131, r_0_132, r_0_133, r_0_134, r_0_135, r_0_136, r_0_137, r_0_138, r_0_139, r_0_140, r_0_141, r_0_142, r_0_143, r_0_144, r_0_145, r_0_146, r_0_147, r_0_148, r_0_149, r_0_150, r_0_151, r_0_152, r_0_153, r_0_154, r_0_155, r_0_156, r_0_157, r_0_158, r_0_159, r_0_160, r_0_161, r_0_162, r_0_163, r_0_164, r_0_165};
  assign row1 = {r_1_0, r_1_1, r_1_2, r_1_3, r_1_4, r_1_5, r_1_6, r_1_7, r_1_8, r_1_9, r_1_10, r_1_11, r_1_12, r_1_13, r_1_14, r_1_15, r_1_16, r_1_17, r_1_18, r_1_19, r_1_20, r_1_21, r_1_22, r_1_23, r_1_24, r_1_25, r_1_26, r_1_27, r_1_28, r_1_29, r_1_30, r_1_31, r_1_32, r_1_33, r_1_34, r_1_35, r_1_36, r_1_37, r_1_38, r_1_39, r_1_40, r_1_41, r_1_42, r_1_43, r_1_44, r_1_45, r_1_46, r_1_47, r_1_48, r_1_49, r_1_50, r_1_51, r_1_52, r_1_53, r_1_54, r_1_55, r_1_56, r_1_57, r_1_58, r_1_59, r_1_60, r_1_61, r_1_62, r_1_63, r_1_64, r_1_65, r_1_66, r_1_67, r_1_68, r_1_69, r_1_70, r_1_71, r_1_72, r_1_73, r_1_74, r_1_75, r_1_76, r_1_77, r_1_78, r_1_79, r_1_80, r_1_81, r_1_82, r_1_83, r_1_84, r_1_85, r_1_86, r_1_87, r_1_88, r_1_89, r_1_90, r_1_91, r_1_92, r_1_93, r_1_94, r_1_95, r_1_96, r_1_97, r_1_98, r_1_99, r_1_100, r_1_101, r_1_102, r_1_103, r_1_104, r_1_105, r_1_106, r_1_107, r_1_108, r_1_109, r_1_110, r_1_111, r_1_112, r_1_113, r_1_114, r_1_115, r_1_116, r_1_117, r_1_118, r_1_119, r_1_120, r_1_121, r_1_122, r_1_123, r_1_124, r_1_125, r_1_126, r_1_127, r_1_128, r_1_129, r_1_130, r_1_131, r_1_132, r_1_133, r_1_134, r_1_135, r_1_136, r_1_137, r_1_138, r_1_139, r_1_140, r_1_141, r_1_142, r_1_143, r_1_144, r_1_145, r_1_146, r_1_147, r_1_148, r_1_149, r_1_150, r_1_151, r_1_152, r_1_153, r_1_154, r_1_155, r_1_156, r_1_157, r_1_158, r_1_159, r_1_160, r_1_161, r_1_162, r_1_163, r_1_164, r_1_165};
  assign row2 = {r_2_0, r_2_1, r_2_2, r_2_3, r_2_4, r_2_5, r_2_6, r_2_7, r_2_8, r_2_9, r_2_10, r_2_11, r_2_12, r_2_13, r_2_14, r_2_15, r_2_16, r_2_17, r_2_18, r_2_19, r_2_20, r_2_21, r_2_22, r_2_23, r_2_24, r_2_25, r_2_26, r_2_27, r_2_28, r_2_29, r_2_30, r_2_31, r_2_32, r_2_33, r_2_34, r_2_35, r_2_36, r_2_37, r_2_38, r_2_39, r_2_40, r_2_41, r_2_42, r_2_43, r_2_44, r_2_45, r_2_46, r_2_47, r_2_48, r_2_49, r_2_50, r_2_51, r_2_52, r_2_53, r_2_54, r_2_55, r_2_56, r_2_57, r_2_58, r_2_59, r_2_60, r_2_61, r_2_62, r_2_63, r_2_64, r_2_65, r_2_66, r_2_67, r_2_68, r_2_69, r_2_70, r_2_71, r_2_72, r_2_73, r_2_74, r_2_75, r_2_76, r_2_77, r_2_78, r_2_79, r_2_80, r_2_81, r_2_82, r_2_83, r_2_84, r_2_85, r_2_86, r_2_87, r_2_88, r_2_89, r_2_90, r_2_91, r_2_92, r_2_93, r_2_94, r_2_95, r_2_96, r_2_97, r_2_98, r_2_99, r_2_100, r_2_101, r_2_102, r_2_103, r_2_104, r_2_105, r_2_106, r_2_107, r_2_108, r_2_109, r_2_110, r_2_111, r_2_112, r_2_113, r_2_114, r_2_115, r_2_116, r_2_117, r_2_118, r_2_119, r_2_120, r_2_121, r_2_122, r_2_123, r_2_124, r_2_125, r_2_126, r_2_127, r_2_128, r_2_129, r_2_130, r_2_131, r_2_132, r_2_133, r_2_134, r_2_135, r_2_136, r_2_137, r_2_138, r_2_139, r_2_140, r_2_141, r_2_142, r_2_143, r_2_144, r_2_145, r_2_146, r_2_147, r_2_148, r_2_149, r_2_150, r_2_151, r_2_152, r_2_153, r_2_154, r_2_155, r_2_156, r_2_157, r_2_158, r_2_159, r_2_160, r_2_161, r_2_162, r_2_163, r_2_164, r_2_165};
  assign row3 = {r_3_0, r_3_1, r_3_2, r_3_3, r_3_4, r_3_5, r_3_6, r_3_7, r_3_8, r_3_9, r_3_10, r_3_11, r_3_12, r_3_13, r_3_14, r_3_15, r_3_16, r_3_17, r_3_18, r_3_19, r_3_20, r_3_21, r_3_22, r_3_23, r_3_24, r_3_25, r_3_26, r_3_27, r_3_28, r_3_29, r_3_30, r_3_31, r_3_32, r_3_33, r_3_34, r_3_35, r_3_36, r_3_37, r_3_38, r_3_39, r_3_40, r_3_41, r_3_42, r_3_43, r_3_44, r_3_45, r_3_46, r_3_47, r_3_48, r_3_49, r_3_50, r_3_51, r_3_52, r_3_53, r_3_54, r_3_55, r_3_56, r_3_57, r_3_58, r_3_59, r_3_60, r_3_61, r_3_62, r_3_63, r_3_64, r_3_65, r_3_66, r_3_67, r_3_68, r_3_69, r_3_70, r_3_71, r_3_72, r_3_73, r_3_74, r_3_75, r_3_76, r_3_77, r_3_78, r_3_79, r_3_80, r_3_81, r_3_82, r_3_83, r_3_84, r_3_85, r_3_86, r_3_87, r_3_88, r_3_89, r_3_90, r_3_91, r_3_92, r_3_93, r_3_94, r_3_95, r_3_96, r_3_97, r_3_98, r_3_99, r_3_100, r_3_101, r_3_102, r_3_103, r_3_104, r_3_105, r_3_106, r_3_107, r_3_108, r_3_109, r_3_110, r_3_111, r_3_112, r_3_113, r_3_114, r_3_115, r_3_116, r_3_117, r_3_118, r_3_119, r_3_120, r_3_121, r_3_122, r_3_123, r_3_124, r_3_125, r_3_126, r_3_127, r_3_128, r_3_129, r_3_130, r_3_131, r_3_132, r_3_133, r_3_134, r_3_135, r_3_136, r_3_137, r_3_138, r_3_139, r_3_140, r_3_141, r_3_142, r_3_143, r_3_144, r_3_145, r_3_146, r_3_147, r_3_148, r_3_149, r_3_150, r_3_151, r_3_152, r_3_153, r_3_154, r_3_155, r_3_156, r_3_157, r_3_158, r_3_159, r_3_160, r_3_161, r_3_162, r_3_163, r_3_164, r_3_165};
  assign row4 = {r_4_0, r_4_1, r_4_2, r_4_3, r_4_4, r_4_5, r_4_6, r_4_7, r_4_8, r_4_9, r_4_10, r_4_11, r_4_12, r_4_13, r_4_14, r_4_15, r_4_16, r_4_17, r_4_18, r_4_19, r_4_20, r_4_21, r_4_22, r_4_23, r_4_24, r_4_25, r_4_26, r_4_27, r_4_28, r_4_29, r_4_30, r_4_31, r_4_32, r_4_33, r_4_34, r_4_35, r_4_36, r_4_37, r_4_38, r_4_39, r_4_40, r_4_41, r_4_42, r_4_43, r_4_44, r_4_45, r_4_46, r_4_47, r_4_48, r_4_49, r_4_50, r_4_51, r_4_52, r_4_53, r_4_54, r_4_55, r_4_56, r_4_57, r_4_58, r_4_59, r_4_60, r_4_61, r_4_62, r_4_63, r_4_64, r_4_65, r_4_66, r_4_67, r_4_68, r_4_69, r_4_70, r_4_71, r_4_72, r_4_73, r_4_74, r_4_75, r_4_76, r_4_77, r_4_78, r_4_79, r_4_80, r_4_81, r_4_82, r_4_83, r_4_84, r_4_85, r_4_86, r_4_87, r_4_88, r_4_89, r_4_90, r_4_91, r_4_92, r_4_93, r_4_94, r_4_95, r_4_96, r_4_97, r_4_98, r_4_99, r_4_100, r_4_101, r_4_102, r_4_103, r_4_104, r_4_105, r_4_106, r_4_107, r_4_108, r_4_109, r_4_110, r_4_111, r_4_112, r_4_113, r_4_114, r_4_115, r_4_116, r_4_117, r_4_118, r_4_119, r_4_120, r_4_121, r_4_122, r_4_123, r_4_124, r_4_125, r_4_126, r_4_127, r_4_128, r_4_129, r_4_130, r_4_131, r_4_132, r_4_133, r_4_134, r_4_135, r_4_136, r_4_137, r_4_138, r_4_139, r_4_140, r_4_141, r_4_142, r_4_143, r_4_144, r_4_145, r_4_146, r_4_147, r_4_148, r_4_149, r_4_150, r_4_151, r_4_152, r_4_153, r_4_154, r_4_155, r_4_156, r_4_157, r_4_158, r_4_159, r_4_160, r_4_161, r_4_162, r_4_163, r_4_164, r_4_165};

  always @(posedge clk) begin
      finish <= ~mode ? start_out_4_165: start_out_0_164;
  end

   //output regular form from skewed form via pipelining
 reg [166:1] result_col0;
 reg [165:1] result_col1;
 reg [164:1] result_col2;
 reg [163:1] result_col3;
 reg [162:1] result_col4;
 reg [161:1] result_col5;
 reg [160:1] result_col6;
 reg [159:1] result_col7;
 reg [158:1] result_col8;
 reg [157:1] result_col9;
 reg [156:1] result_col10;
 reg [155:1] result_col11;
 reg [154:1] result_col12;
 reg [153:1] result_col13;
 reg [152:1] result_col14;
 reg [151:1] result_col15;
 reg [150:1] result_col16;
 reg [149:1] result_col17;
 reg [148:1] result_col18;
 reg [147:1] result_col19;
 reg [146:1] result_col20;
 reg [145:1] result_col21;
 reg [144:1] result_col22;
 reg [143:1] result_col23;
 reg [142:1] result_col24;
 reg [141:1] result_col25;
 reg [140:1] result_col26;
 reg [139:1] result_col27;
 reg [138:1] result_col28;
 reg [137:1] result_col29;
 reg [136:1] result_col30;
 reg [135:1] result_col31;
 reg [134:1] result_col32;
 reg [133:1] result_col33;
 reg [132:1] result_col34;
 reg [131:1] result_col35;
 reg [130:1] result_col36;
 reg [129:1] result_col37;
 reg [128:1] result_col38;
 reg [127:1] result_col39;
 reg [126:1] result_col40;
 reg [125:1] result_col41;
 reg [124:1] result_col42;
 reg [123:1] result_col43;
 reg [122:1] result_col44;
 reg [121:1] result_col45;
 reg [120:1] result_col46;
 reg [119:1] result_col47;
 reg [118:1] result_col48;
 reg [117:1] result_col49;
 reg [116:1] result_col50;
 reg [115:1] result_col51;
 reg [114:1] result_col52;
 reg [113:1] result_col53;
 reg [112:1] result_col54;
 reg [111:1] result_col55;
 reg [110:1] result_col56;
 reg [109:1] result_col57;
 reg [108:1] result_col58;
 reg [107:1] result_col59;
 reg [106:1] result_col60;
 reg [105:1] result_col61;
 reg [104:1] result_col62;
 reg [103:1] result_col63;
 reg [102:1] result_col64;
 reg [101:1] result_col65;
 reg [100:1] result_col66;
 reg [99:1] result_col67;
 reg [98:1] result_col68;
 reg [97:1] result_col69;
 reg [96:1] result_col70;
 reg [95:1] result_col71;
 reg [94:1] result_col72;
 reg [93:1] result_col73;
 reg [92:1] result_col74;
 reg [91:1] result_col75;
 reg [90:1] result_col76;
 reg [89:1] result_col77;
 reg [88:1] result_col78;
 reg [87:1] result_col79;
 reg [86:1] result_col80;
 reg [85:1] result_col81;
 reg [84:1] result_col82;
 reg [83:1] result_col83;
 reg [82:1] result_col84;
 reg [81:1] result_col85;
 reg [80:1] result_col86;
 reg [79:1] result_col87;
 reg [78:1] result_col88;
 reg [77:1] result_col89;
 reg [76:1] result_col90;
 reg [75:1] result_col91;
 reg [74:1] result_col92;
 reg [73:1] result_col93;
 reg [72:1] result_col94;
 reg [71:1] result_col95;
 reg [70:1] result_col96;
 reg [69:1] result_col97;
 reg [68:1] result_col98;
 reg [67:1] result_col99;
 reg [66:1] result_col100;
 reg [65:1] result_col101;
 reg [64:1] result_col102;
 reg [63:1] result_col103;
 reg [62:1] result_col104;
 reg [61:1] result_col105;
 reg [60:1] result_col106;
 reg [59:1] result_col107;
 reg [58:1] result_col108;
 reg [57:1] result_col109;
 reg [56:1] result_col110;
 reg [55:1] result_col111;
 reg [54:1] result_col112;
 reg [53:1] result_col113;
 reg [52:1] result_col114;
 reg [51:1] result_col115;
 reg [50:1] result_col116;
 reg [49:1] result_col117;
 reg [48:1] result_col118;
 reg [47:1] result_col119;
 reg [46:1] result_col120;
 reg [45:1] result_col121;
 reg [44:1] result_col122;
 reg [43:1] result_col123;
 reg [42:1] result_col124;
 reg [41:1] result_col125;
 reg [40:1] result_col126;
 reg [39:1] result_col127;
 reg [38:1] result_col128;
 reg [37:1] result_col129;
 reg [36:1] result_col130;
 reg [35:1] result_col131;
 reg [34:1] result_col132;
 reg [33:1] result_col133;
 reg [32:1] result_col134;
 reg [31:1] result_col135;
 reg [30:1] result_col136;
 reg [29:1] result_col137;
 reg [28:1] result_col138;
 reg [27:1] result_col139;
 reg [26:1] result_col140;
 reg [25:1] result_col141;
 reg [24:1] result_col142;
 reg [23:1] result_col143;
 reg [22:1] result_col144;
 reg [21:1] result_col145;
 reg [20:1] result_col146;
 reg [19:1] result_col147;
 reg [18:1] result_col148;
 reg [17:1] result_col149;
 reg [16:1] result_col150;
 reg [15:1] result_col151;
 reg [14:1] result_col152;
 reg [13:1] result_col153;
 reg [12:1] result_col154;
 reg [11:1] result_col155;
 reg [10:1] result_col156;
 reg [9:1] result_col157;
 reg [8:1] result_col158;
 reg [7:1] result_col159;
 reg [6:1] result_col160;
 reg [5:1] result_col161;
 reg [4:1] result_col162;
 reg [3:1] result_col163;
 reg [2:1] result_col164;
 reg [1:1] result_col165;

  always @(posedge clk) begin
   result_col0[1] <= data_out_4_0;
   result_col0[2] <= result_col0[1];
   result_col0[3] <= result_col0[2];
   result_col0[4] <= result_col0[3];
   result_col0[5] <= result_col0[4];
   result_col0[6] <= result_col0[5];
   result_col0[7] <= result_col0[6];
   result_col0[8] <= result_col0[7];
   result_col0[9] <= result_col0[8];
   result_col0[10] <= result_col0[9];
   result_col0[11] <= result_col0[10];
   result_col0[12] <= result_col0[11];
   result_col0[13] <= result_col0[12];
   result_col0[14] <= result_col0[13];
   result_col0[15] <= result_col0[14];
   result_col0[16] <= result_col0[15];
   result_col0[17] <= result_col0[16];
   result_col0[18] <= result_col0[17];
   result_col0[19] <= result_col0[18];
   result_col0[20] <= result_col0[19];
   result_col0[21] <= result_col0[20];
   result_col0[22] <= result_col0[21];
   result_col0[23] <= result_col0[22];
   result_col0[24] <= result_col0[23];
   result_col0[25] <= result_col0[24];
   result_col0[26] <= result_col0[25];
   result_col0[27] <= result_col0[26];
   result_col0[28] <= result_col0[27];
   result_col0[29] <= result_col0[28];
   result_col0[30] <= result_col0[29];
   result_col0[31] <= result_col0[30];
   result_col0[32] <= result_col0[31];
   result_col0[33] <= result_col0[32];
   result_col0[34] <= result_col0[33];
   result_col0[35] <= result_col0[34];
   result_col0[36] <= result_col0[35];
   result_col0[37] <= result_col0[36];
   result_col0[38] <= result_col0[37];
   result_col0[39] <= result_col0[38];
   result_col0[40] <= result_col0[39];
   result_col0[41] <= result_col0[40];
   result_col0[42] <= result_col0[41];
   result_col0[43] <= result_col0[42];
   result_col0[44] <= result_col0[43];
   result_col0[45] <= result_col0[44];
   result_col0[46] <= result_col0[45];
   result_col0[47] <= result_col0[46];
   result_col0[48] <= result_col0[47];
   result_col0[49] <= result_col0[48];
   result_col0[50] <= result_col0[49];
   result_col0[51] <= result_col0[50];
   result_col0[52] <= result_col0[51];
   result_col0[53] <= result_col0[52];
   result_col0[54] <= result_col0[53];
   result_col0[55] <= result_col0[54];
   result_col0[56] <= result_col0[55];
   result_col0[57] <= result_col0[56];
   result_col0[58] <= result_col0[57];
   result_col0[59] <= result_col0[58];
   result_col0[60] <= result_col0[59];
   result_col0[61] <= result_col0[60];
   result_col0[62] <= result_col0[61];
   result_col0[63] <= result_col0[62];
   result_col0[64] <= result_col0[63];
   result_col0[65] <= result_col0[64];
   result_col0[66] <= result_col0[65];
   result_col0[67] <= result_col0[66];
   result_col0[68] <= result_col0[67];
   result_col0[69] <= result_col0[68];
   result_col0[70] <= result_col0[69];
   result_col0[71] <= result_col0[70];
   result_col0[72] <= result_col0[71];
   result_col0[73] <= result_col0[72];
   result_col0[74] <= result_col0[73];
   result_col0[75] <= result_col0[74];
   result_col0[76] <= result_col0[75];
   result_col0[77] <= result_col0[76];
   result_col0[78] <= result_col0[77];
   result_col0[79] <= result_col0[78];
   result_col0[80] <= result_col0[79];
   result_col0[81] <= result_col0[80];
   result_col0[82] <= result_col0[81];
   result_col0[83] <= result_col0[82];
   result_col0[84] <= result_col0[83];
   result_col0[85] <= result_col0[84];
   result_col0[86] <= result_col0[85];
   result_col0[87] <= result_col0[86];
   result_col0[88] <= result_col0[87];
   result_col0[89] <= result_col0[88];
   result_col0[90] <= result_col0[89];
   result_col0[91] <= result_col0[90];
   result_col0[92] <= result_col0[91];
   result_col0[93] <= result_col0[92];
   result_col0[94] <= result_col0[93];
   result_col0[95] <= result_col0[94];
   result_col0[96] <= result_col0[95];
   result_col0[97] <= result_col0[96];
   result_col0[98] <= result_col0[97];
   result_col0[99] <= result_col0[98];
   result_col0[100] <= result_col0[99];
   result_col0[101] <= result_col0[100];
   result_col0[102] <= result_col0[101];
   result_col0[103] <= result_col0[102];
   result_col0[104] <= result_col0[103];
   result_col0[105] <= result_col0[104];
   result_col0[106] <= result_col0[105];
   result_col0[107] <= result_col0[106];
   result_col0[108] <= result_col0[107];
   result_col0[109] <= result_col0[108];
   result_col0[110] <= result_col0[109];
   result_col0[111] <= result_col0[110];
   result_col0[112] <= result_col0[111];
   result_col0[113] <= result_col0[112];
   result_col0[114] <= result_col0[113];
   result_col0[115] <= result_col0[114];
   result_col0[116] <= result_col0[115];
   result_col0[117] <= result_col0[116];
   result_col0[118] <= result_col0[117];
   result_col0[119] <= result_col0[118];
   result_col0[120] <= result_col0[119];
   result_col0[121] <= result_col0[120];
   result_col0[122] <= result_col0[121];
   result_col0[123] <= result_col0[122];
   result_col0[124] <= result_col0[123];
   result_col0[125] <= result_col0[124];
   result_col0[126] <= result_col0[125];
   result_col0[127] <= result_col0[126];
   result_col0[128] <= result_col0[127];
   result_col0[129] <= result_col0[128];
   result_col0[130] <= result_col0[129];
   result_col0[131] <= result_col0[130];
   result_col0[132] <= result_col0[131];
   result_col0[133] <= result_col0[132];
   result_col0[134] <= result_col0[133];
   result_col0[135] <= result_col0[134];
   result_col0[136] <= result_col0[135];
   result_col0[137] <= result_col0[136];
   result_col0[138] <= result_col0[137];
   result_col0[139] <= result_col0[138];
   result_col0[140] <= result_col0[139];
   result_col0[141] <= result_col0[140];
   result_col0[142] <= result_col0[141];
   result_col0[143] <= result_col0[142];
   result_col0[144] <= result_col0[143];
   result_col0[145] <= result_col0[144];
   result_col0[146] <= result_col0[145];
   result_col0[147] <= result_col0[146];
   result_col0[148] <= result_col0[147];
   result_col0[149] <= result_col0[148];
   result_col0[150] <= result_col0[149];
   result_col0[151] <= result_col0[150];
   result_col0[152] <= result_col0[151];
   result_col0[153] <= result_col0[152];
   result_col0[154] <= result_col0[153];
   result_col0[155] <= result_col0[154];
   result_col0[156] <= result_col0[155];
   result_col0[157] <= result_col0[156];
   result_col0[158] <= result_col0[157];
   result_col0[159] <= result_col0[158];
   result_col0[160] <= result_col0[159];
   result_col0[161] <= result_col0[160];
   result_col0[162] <= result_col0[161];
   result_col0[163] <= result_col0[162];
   result_col0[164] <= result_col0[163];
   result_col0[165] <= result_col0[164];
   result_col0[166] <= result_col0[165];

   result_col1[1] <= data_out_4_1;
   result_col1[2] <= result_col1[1];
   result_col1[3] <= result_col1[2];
   result_col1[4] <= result_col1[3];
   result_col1[5] <= result_col1[4];
   result_col1[6] <= result_col1[5];
   result_col1[7] <= result_col1[6];
   result_col1[8] <= result_col1[7];
   result_col1[9] <= result_col1[8];
   result_col1[10] <= result_col1[9];
   result_col1[11] <= result_col1[10];
   result_col1[12] <= result_col1[11];
   result_col1[13] <= result_col1[12];
   result_col1[14] <= result_col1[13];
   result_col1[15] <= result_col1[14];
   result_col1[16] <= result_col1[15];
   result_col1[17] <= result_col1[16];
   result_col1[18] <= result_col1[17];
   result_col1[19] <= result_col1[18];
   result_col1[20] <= result_col1[19];
   result_col1[21] <= result_col1[20];
   result_col1[22] <= result_col1[21];
   result_col1[23] <= result_col1[22];
   result_col1[24] <= result_col1[23];
   result_col1[25] <= result_col1[24];
   result_col1[26] <= result_col1[25];
   result_col1[27] <= result_col1[26];
   result_col1[28] <= result_col1[27];
   result_col1[29] <= result_col1[28];
   result_col1[30] <= result_col1[29];
   result_col1[31] <= result_col1[30];
   result_col1[32] <= result_col1[31];
   result_col1[33] <= result_col1[32];
   result_col1[34] <= result_col1[33];
   result_col1[35] <= result_col1[34];
   result_col1[36] <= result_col1[35];
   result_col1[37] <= result_col1[36];
   result_col1[38] <= result_col1[37];
   result_col1[39] <= result_col1[38];
   result_col1[40] <= result_col1[39];
   result_col1[41] <= result_col1[40];
   result_col1[42] <= result_col1[41];
   result_col1[43] <= result_col1[42];
   result_col1[44] <= result_col1[43];
   result_col1[45] <= result_col1[44];
   result_col1[46] <= result_col1[45];
   result_col1[47] <= result_col1[46];
   result_col1[48] <= result_col1[47];
   result_col1[49] <= result_col1[48];
   result_col1[50] <= result_col1[49];
   result_col1[51] <= result_col1[50];
   result_col1[52] <= result_col1[51];
   result_col1[53] <= result_col1[52];
   result_col1[54] <= result_col1[53];
   result_col1[55] <= result_col1[54];
   result_col1[56] <= result_col1[55];
   result_col1[57] <= result_col1[56];
   result_col1[58] <= result_col1[57];
   result_col1[59] <= result_col1[58];
   result_col1[60] <= result_col1[59];
   result_col1[61] <= result_col1[60];
   result_col1[62] <= result_col1[61];
   result_col1[63] <= result_col1[62];
   result_col1[64] <= result_col1[63];
   result_col1[65] <= result_col1[64];
   result_col1[66] <= result_col1[65];
   result_col1[67] <= result_col1[66];
   result_col1[68] <= result_col1[67];
   result_col1[69] <= result_col1[68];
   result_col1[70] <= result_col1[69];
   result_col1[71] <= result_col1[70];
   result_col1[72] <= result_col1[71];
   result_col1[73] <= result_col1[72];
   result_col1[74] <= result_col1[73];
   result_col1[75] <= result_col1[74];
   result_col1[76] <= result_col1[75];
   result_col1[77] <= result_col1[76];
   result_col1[78] <= result_col1[77];
   result_col1[79] <= result_col1[78];
   result_col1[80] <= result_col1[79];
   result_col1[81] <= result_col1[80];
   result_col1[82] <= result_col1[81];
   result_col1[83] <= result_col1[82];
   result_col1[84] <= result_col1[83];
   result_col1[85] <= result_col1[84];
   result_col1[86] <= result_col1[85];
   result_col1[87] <= result_col1[86];
   result_col1[88] <= result_col1[87];
   result_col1[89] <= result_col1[88];
   result_col1[90] <= result_col1[89];
   result_col1[91] <= result_col1[90];
   result_col1[92] <= result_col1[91];
   result_col1[93] <= result_col1[92];
   result_col1[94] <= result_col1[93];
   result_col1[95] <= result_col1[94];
   result_col1[96] <= result_col1[95];
   result_col1[97] <= result_col1[96];
   result_col1[98] <= result_col1[97];
   result_col1[99] <= result_col1[98];
   result_col1[100] <= result_col1[99];
   result_col1[101] <= result_col1[100];
   result_col1[102] <= result_col1[101];
   result_col1[103] <= result_col1[102];
   result_col1[104] <= result_col1[103];
   result_col1[105] <= result_col1[104];
   result_col1[106] <= result_col1[105];
   result_col1[107] <= result_col1[106];
   result_col1[108] <= result_col1[107];
   result_col1[109] <= result_col1[108];
   result_col1[110] <= result_col1[109];
   result_col1[111] <= result_col1[110];
   result_col1[112] <= result_col1[111];
   result_col1[113] <= result_col1[112];
   result_col1[114] <= result_col1[113];
   result_col1[115] <= result_col1[114];
   result_col1[116] <= result_col1[115];
   result_col1[117] <= result_col1[116];
   result_col1[118] <= result_col1[117];
   result_col1[119] <= result_col1[118];
   result_col1[120] <= result_col1[119];
   result_col1[121] <= result_col1[120];
   result_col1[122] <= result_col1[121];
   result_col1[123] <= result_col1[122];
   result_col1[124] <= result_col1[123];
   result_col1[125] <= result_col1[124];
   result_col1[126] <= result_col1[125];
   result_col1[127] <= result_col1[126];
   result_col1[128] <= result_col1[127];
   result_col1[129] <= result_col1[128];
   result_col1[130] <= result_col1[129];
   result_col1[131] <= result_col1[130];
   result_col1[132] <= result_col1[131];
   result_col1[133] <= result_col1[132];
   result_col1[134] <= result_col1[133];
   result_col1[135] <= result_col1[134];
   result_col1[136] <= result_col1[135];
   result_col1[137] <= result_col1[136];
   result_col1[138] <= result_col1[137];
   result_col1[139] <= result_col1[138];
   result_col1[140] <= result_col1[139];
   result_col1[141] <= result_col1[140];
   result_col1[142] <= result_col1[141];
   result_col1[143] <= result_col1[142];
   result_col1[144] <= result_col1[143];
   result_col1[145] <= result_col1[144];
   result_col1[146] <= result_col1[145];
   result_col1[147] <= result_col1[146];
   result_col1[148] <= result_col1[147];
   result_col1[149] <= result_col1[148];
   result_col1[150] <= result_col1[149];
   result_col1[151] <= result_col1[150];
   result_col1[152] <= result_col1[151];
   result_col1[153] <= result_col1[152];
   result_col1[154] <= result_col1[153];
   result_col1[155] <= result_col1[154];
   result_col1[156] <= result_col1[155];
   result_col1[157] <= result_col1[156];
   result_col1[158] <= result_col1[157];
   result_col1[159] <= result_col1[158];
   result_col1[160] <= result_col1[159];
   result_col1[161] <= result_col1[160];
   result_col1[162] <= result_col1[161];
   result_col1[163] <= result_col1[162];
   result_col1[164] <= result_col1[163];
   result_col1[165] <= result_col1[164];

   result_col2[1] <= data_out_4_2;
   result_col2[2] <= result_col2[1];
   result_col2[3] <= result_col2[2];
   result_col2[4] <= result_col2[3];
   result_col2[5] <= result_col2[4];
   result_col2[6] <= result_col2[5];
   result_col2[7] <= result_col2[6];
   result_col2[8] <= result_col2[7];
   result_col2[9] <= result_col2[8];
   result_col2[10] <= result_col2[9];
   result_col2[11] <= result_col2[10];
   result_col2[12] <= result_col2[11];
   result_col2[13] <= result_col2[12];
   result_col2[14] <= result_col2[13];
   result_col2[15] <= result_col2[14];
   result_col2[16] <= result_col2[15];
   result_col2[17] <= result_col2[16];
   result_col2[18] <= result_col2[17];
   result_col2[19] <= result_col2[18];
   result_col2[20] <= result_col2[19];
   result_col2[21] <= result_col2[20];
   result_col2[22] <= result_col2[21];
   result_col2[23] <= result_col2[22];
   result_col2[24] <= result_col2[23];
   result_col2[25] <= result_col2[24];
   result_col2[26] <= result_col2[25];
   result_col2[27] <= result_col2[26];
   result_col2[28] <= result_col2[27];
   result_col2[29] <= result_col2[28];
   result_col2[30] <= result_col2[29];
   result_col2[31] <= result_col2[30];
   result_col2[32] <= result_col2[31];
   result_col2[33] <= result_col2[32];
   result_col2[34] <= result_col2[33];
   result_col2[35] <= result_col2[34];
   result_col2[36] <= result_col2[35];
   result_col2[37] <= result_col2[36];
   result_col2[38] <= result_col2[37];
   result_col2[39] <= result_col2[38];
   result_col2[40] <= result_col2[39];
   result_col2[41] <= result_col2[40];
   result_col2[42] <= result_col2[41];
   result_col2[43] <= result_col2[42];
   result_col2[44] <= result_col2[43];
   result_col2[45] <= result_col2[44];
   result_col2[46] <= result_col2[45];
   result_col2[47] <= result_col2[46];
   result_col2[48] <= result_col2[47];
   result_col2[49] <= result_col2[48];
   result_col2[50] <= result_col2[49];
   result_col2[51] <= result_col2[50];
   result_col2[52] <= result_col2[51];
   result_col2[53] <= result_col2[52];
   result_col2[54] <= result_col2[53];
   result_col2[55] <= result_col2[54];
   result_col2[56] <= result_col2[55];
   result_col2[57] <= result_col2[56];
   result_col2[58] <= result_col2[57];
   result_col2[59] <= result_col2[58];
   result_col2[60] <= result_col2[59];
   result_col2[61] <= result_col2[60];
   result_col2[62] <= result_col2[61];
   result_col2[63] <= result_col2[62];
   result_col2[64] <= result_col2[63];
   result_col2[65] <= result_col2[64];
   result_col2[66] <= result_col2[65];
   result_col2[67] <= result_col2[66];
   result_col2[68] <= result_col2[67];
   result_col2[69] <= result_col2[68];
   result_col2[70] <= result_col2[69];
   result_col2[71] <= result_col2[70];
   result_col2[72] <= result_col2[71];
   result_col2[73] <= result_col2[72];
   result_col2[74] <= result_col2[73];
   result_col2[75] <= result_col2[74];
   result_col2[76] <= result_col2[75];
   result_col2[77] <= result_col2[76];
   result_col2[78] <= result_col2[77];
   result_col2[79] <= result_col2[78];
   result_col2[80] <= result_col2[79];
   result_col2[81] <= result_col2[80];
   result_col2[82] <= result_col2[81];
   result_col2[83] <= result_col2[82];
   result_col2[84] <= result_col2[83];
   result_col2[85] <= result_col2[84];
   result_col2[86] <= result_col2[85];
   result_col2[87] <= result_col2[86];
   result_col2[88] <= result_col2[87];
   result_col2[89] <= result_col2[88];
   result_col2[90] <= result_col2[89];
   result_col2[91] <= result_col2[90];
   result_col2[92] <= result_col2[91];
   result_col2[93] <= result_col2[92];
   result_col2[94] <= result_col2[93];
   result_col2[95] <= result_col2[94];
   result_col2[96] <= result_col2[95];
   result_col2[97] <= result_col2[96];
   result_col2[98] <= result_col2[97];
   result_col2[99] <= result_col2[98];
   result_col2[100] <= result_col2[99];
   result_col2[101] <= result_col2[100];
   result_col2[102] <= result_col2[101];
   result_col2[103] <= result_col2[102];
   result_col2[104] <= result_col2[103];
   result_col2[105] <= result_col2[104];
   result_col2[106] <= result_col2[105];
   result_col2[107] <= result_col2[106];
   result_col2[108] <= result_col2[107];
   result_col2[109] <= result_col2[108];
   result_col2[110] <= result_col2[109];
   result_col2[111] <= result_col2[110];
   result_col2[112] <= result_col2[111];
   result_col2[113] <= result_col2[112];
   result_col2[114] <= result_col2[113];
   result_col2[115] <= result_col2[114];
   result_col2[116] <= result_col2[115];
   result_col2[117] <= result_col2[116];
   result_col2[118] <= result_col2[117];
   result_col2[119] <= result_col2[118];
   result_col2[120] <= result_col2[119];
   result_col2[121] <= result_col2[120];
   result_col2[122] <= result_col2[121];
   result_col2[123] <= result_col2[122];
   result_col2[124] <= result_col2[123];
   result_col2[125] <= result_col2[124];
   result_col2[126] <= result_col2[125];
   result_col2[127] <= result_col2[126];
   result_col2[128] <= result_col2[127];
   result_col2[129] <= result_col2[128];
   result_col2[130] <= result_col2[129];
   result_col2[131] <= result_col2[130];
   result_col2[132] <= result_col2[131];
   result_col2[133] <= result_col2[132];
   result_col2[134] <= result_col2[133];
   result_col2[135] <= result_col2[134];
   result_col2[136] <= result_col2[135];
   result_col2[137] <= result_col2[136];
   result_col2[138] <= result_col2[137];
   result_col2[139] <= result_col2[138];
   result_col2[140] <= result_col2[139];
   result_col2[141] <= result_col2[140];
   result_col2[142] <= result_col2[141];
   result_col2[143] <= result_col2[142];
   result_col2[144] <= result_col2[143];
   result_col2[145] <= result_col2[144];
   result_col2[146] <= result_col2[145];
   result_col2[147] <= result_col2[146];
   result_col2[148] <= result_col2[147];
   result_col2[149] <= result_col2[148];
   result_col2[150] <= result_col2[149];
   result_col2[151] <= result_col2[150];
   result_col2[152] <= result_col2[151];
   result_col2[153] <= result_col2[152];
   result_col2[154] <= result_col2[153];
   result_col2[155] <= result_col2[154];
   result_col2[156] <= result_col2[155];
   result_col2[157] <= result_col2[156];
   result_col2[158] <= result_col2[157];
   result_col2[159] <= result_col2[158];
   result_col2[160] <= result_col2[159];
   result_col2[161] <= result_col2[160];
   result_col2[162] <= result_col2[161];
   result_col2[163] <= result_col2[162];
   result_col2[164] <= result_col2[163];

   result_col3[1] <= data_out_4_3;
   result_col3[2] <= result_col3[1];
   result_col3[3] <= result_col3[2];
   result_col3[4] <= result_col3[3];
   result_col3[5] <= result_col3[4];
   result_col3[6] <= result_col3[5];
   result_col3[7] <= result_col3[6];
   result_col3[8] <= result_col3[7];
   result_col3[9] <= result_col3[8];
   result_col3[10] <= result_col3[9];
   result_col3[11] <= result_col3[10];
   result_col3[12] <= result_col3[11];
   result_col3[13] <= result_col3[12];
   result_col3[14] <= result_col3[13];
   result_col3[15] <= result_col3[14];
   result_col3[16] <= result_col3[15];
   result_col3[17] <= result_col3[16];
   result_col3[18] <= result_col3[17];
   result_col3[19] <= result_col3[18];
   result_col3[20] <= result_col3[19];
   result_col3[21] <= result_col3[20];
   result_col3[22] <= result_col3[21];
   result_col3[23] <= result_col3[22];
   result_col3[24] <= result_col3[23];
   result_col3[25] <= result_col3[24];
   result_col3[26] <= result_col3[25];
   result_col3[27] <= result_col3[26];
   result_col3[28] <= result_col3[27];
   result_col3[29] <= result_col3[28];
   result_col3[30] <= result_col3[29];
   result_col3[31] <= result_col3[30];
   result_col3[32] <= result_col3[31];
   result_col3[33] <= result_col3[32];
   result_col3[34] <= result_col3[33];
   result_col3[35] <= result_col3[34];
   result_col3[36] <= result_col3[35];
   result_col3[37] <= result_col3[36];
   result_col3[38] <= result_col3[37];
   result_col3[39] <= result_col3[38];
   result_col3[40] <= result_col3[39];
   result_col3[41] <= result_col3[40];
   result_col3[42] <= result_col3[41];
   result_col3[43] <= result_col3[42];
   result_col3[44] <= result_col3[43];
   result_col3[45] <= result_col3[44];
   result_col3[46] <= result_col3[45];
   result_col3[47] <= result_col3[46];
   result_col3[48] <= result_col3[47];
   result_col3[49] <= result_col3[48];
   result_col3[50] <= result_col3[49];
   result_col3[51] <= result_col3[50];
   result_col3[52] <= result_col3[51];
   result_col3[53] <= result_col3[52];
   result_col3[54] <= result_col3[53];
   result_col3[55] <= result_col3[54];
   result_col3[56] <= result_col3[55];
   result_col3[57] <= result_col3[56];
   result_col3[58] <= result_col3[57];
   result_col3[59] <= result_col3[58];
   result_col3[60] <= result_col3[59];
   result_col3[61] <= result_col3[60];
   result_col3[62] <= result_col3[61];
   result_col3[63] <= result_col3[62];
   result_col3[64] <= result_col3[63];
   result_col3[65] <= result_col3[64];
   result_col3[66] <= result_col3[65];
   result_col3[67] <= result_col3[66];
   result_col3[68] <= result_col3[67];
   result_col3[69] <= result_col3[68];
   result_col3[70] <= result_col3[69];
   result_col3[71] <= result_col3[70];
   result_col3[72] <= result_col3[71];
   result_col3[73] <= result_col3[72];
   result_col3[74] <= result_col3[73];
   result_col3[75] <= result_col3[74];
   result_col3[76] <= result_col3[75];
   result_col3[77] <= result_col3[76];
   result_col3[78] <= result_col3[77];
   result_col3[79] <= result_col3[78];
   result_col3[80] <= result_col3[79];
   result_col3[81] <= result_col3[80];
   result_col3[82] <= result_col3[81];
   result_col3[83] <= result_col3[82];
   result_col3[84] <= result_col3[83];
   result_col3[85] <= result_col3[84];
   result_col3[86] <= result_col3[85];
   result_col3[87] <= result_col3[86];
   result_col3[88] <= result_col3[87];
   result_col3[89] <= result_col3[88];
   result_col3[90] <= result_col3[89];
   result_col3[91] <= result_col3[90];
   result_col3[92] <= result_col3[91];
   result_col3[93] <= result_col3[92];
   result_col3[94] <= result_col3[93];
   result_col3[95] <= result_col3[94];
   result_col3[96] <= result_col3[95];
   result_col3[97] <= result_col3[96];
   result_col3[98] <= result_col3[97];
   result_col3[99] <= result_col3[98];
   result_col3[100] <= result_col3[99];
   result_col3[101] <= result_col3[100];
   result_col3[102] <= result_col3[101];
   result_col3[103] <= result_col3[102];
   result_col3[104] <= result_col3[103];
   result_col3[105] <= result_col3[104];
   result_col3[106] <= result_col3[105];
   result_col3[107] <= result_col3[106];
   result_col3[108] <= result_col3[107];
   result_col3[109] <= result_col3[108];
   result_col3[110] <= result_col3[109];
   result_col3[111] <= result_col3[110];
   result_col3[112] <= result_col3[111];
   result_col3[113] <= result_col3[112];
   result_col3[114] <= result_col3[113];
   result_col3[115] <= result_col3[114];
   result_col3[116] <= result_col3[115];
   result_col3[117] <= result_col3[116];
   result_col3[118] <= result_col3[117];
   result_col3[119] <= result_col3[118];
   result_col3[120] <= result_col3[119];
   result_col3[121] <= result_col3[120];
   result_col3[122] <= result_col3[121];
   result_col3[123] <= result_col3[122];
   result_col3[124] <= result_col3[123];
   result_col3[125] <= result_col3[124];
   result_col3[126] <= result_col3[125];
   result_col3[127] <= result_col3[126];
   result_col3[128] <= result_col3[127];
   result_col3[129] <= result_col3[128];
   result_col3[130] <= result_col3[129];
   result_col3[131] <= result_col3[130];
   result_col3[132] <= result_col3[131];
   result_col3[133] <= result_col3[132];
   result_col3[134] <= result_col3[133];
   result_col3[135] <= result_col3[134];
   result_col3[136] <= result_col3[135];
   result_col3[137] <= result_col3[136];
   result_col3[138] <= result_col3[137];
   result_col3[139] <= result_col3[138];
   result_col3[140] <= result_col3[139];
   result_col3[141] <= result_col3[140];
   result_col3[142] <= result_col3[141];
   result_col3[143] <= result_col3[142];
   result_col3[144] <= result_col3[143];
   result_col3[145] <= result_col3[144];
   result_col3[146] <= result_col3[145];
   result_col3[147] <= result_col3[146];
   result_col3[148] <= result_col3[147];
   result_col3[149] <= result_col3[148];
   result_col3[150] <= result_col3[149];
   result_col3[151] <= result_col3[150];
   result_col3[152] <= result_col3[151];
   result_col3[153] <= result_col3[152];
   result_col3[154] <= result_col3[153];
   result_col3[155] <= result_col3[154];
   result_col3[156] <= result_col3[155];
   result_col3[157] <= result_col3[156];
   result_col3[158] <= result_col3[157];
   result_col3[159] <= result_col3[158];
   result_col3[160] <= result_col3[159];
   result_col3[161] <= result_col3[160];
   result_col3[162] <= result_col3[161];
   result_col3[163] <= result_col3[162];

   result_col4[1] <= data_out_4_4;
   result_col4[2] <= result_col4[1];
   result_col4[3] <= result_col4[2];
   result_col4[4] <= result_col4[3];
   result_col4[5] <= result_col4[4];
   result_col4[6] <= result_col4[5];
   result_col4[7] <= result_col4[6];
   result_col4[8] <= result_col4[7];
   result_col4[9] <= result_col4[8];
   result_col4[10] <= result_col4[9];
   result_col4[11] <= result_col4[10];
   result_col4[12] <= result_col4[11];
   result_col4[13] <= result_col4[12];
   result_col4[14] <= result_col4[13];
   result_col4[15] <= result_col4[14];
   result_col4[16] <= result_col4[15];
   result_col4[17] <= result_col4[16];
   result_col4[18] <= result_col4[17];
   result_col4[19] <= result_col4[18];
   result_col4[20] <= result_col4[19];
   result_col4[21] <= result_col4[20];
   result_col4[22] <= result_col4[21];
   result_col4[23] <= result_col4[22];
   result_col4[24] <= result_col4[23];
   result_col4[25] <= result_col4[24];
   result_col4[26] <= result_col4[25];
   result_col4[27] <= result_col4[26];
   result_col4[28] <= result_col4[27];
   result_col4[29] <= result_col4[28];
   result_col4[30] <= result_col4[29];
   result_col4[31] <= result_col4[30];
   result_col4[32] <= result_col4[31];
   result_col4[33] <= result_col4[32];
   result_col4[34] <= result_col4[33];
   result_col4[35] <= result_col4[34];
   result_col4[36] <= result_col4[35];
   result_col4[37] <= result_col4[36];
   result_col4[38] <= result_col4[37];
   result_col4[39] <= result_col4[38];
   result_col4[40] <= result_col4[39];
   result_col4[41] <= result_col4[40];
   result_col4[42] <= result_col4[41];
   result_col4[43] <= result_col4[42];
   result_col4[44] <= result_col4[43];
   result_col4[45] <= result_col4[44];
   result_col4[46] <= result_col4[45];
   result_col4[47] <= result_col4[46];
   result_col4[48] <= result_col4[47];
   result_col4[49] <= result_col4[48];
   result_col4[50] <= result_col4[49];
   result_col4[51] <= result_col4[50];
   result_col4[52] <= result_col4[51];
   result_col4[53] <= result_col4[52];
   result_col4[54] <= result_col4[53];
   result_col4[55] <= result_col4[54];
   result_col4[56] <= result_col4[55];
   result_col4[57] <= result_col4[56];
   result_col4[58] <= result_col4[57];
   result_col4[59] <= result_col4[58];
   result_col4[60] <= result_col4[59];
   result_col4[61] <= result_col4[60];
   result_col4[62] <= result_col4[61];
   result_col4[63] <= result_col4[62];
   result_col4[64] <= result_col4[63];
   result_col4[65] <= result_col4[64];
   result_col4[66] <= result_col4[65];
   result_col4[67] <= result_col4[66];
   result_col4[68] <= result_col4[67];
   result_col4[69] <= result_col4[68];
   result_col4[70] <= result_col4[69];
   result_col4[71] <= result_col4[70];
   result_col4[72] <= result_col4[71];
   result_col4[73] <= result_col4[72];
   result_col4[74] <= result_col4[73];
   result_col4[75] <= result_col4[74];
   result_col4[76] <= result_col4[75];
   result_col4[77] <= result_col4[76];
   result_col4[78] <= result_col4[77];
   result_col4[79] <= result_col4[78];
   result_col4[80] <= result_col4[79];
   result_col4[81] <= result_col4[80];
   result_col4[82] <= result_col4[81];
   result_col4[83] <= result_col4[82];
   result_col4[84] <= result_col4[83];
   result_col4[85] <= result_col4[84];
   result_col4[86] <= result_col4[85];
   result_col4[87] <= result_col4[86];
   result_col4[88] <= result_col4[87];
   result_col4[89] <= result_col4[88];
   result_col4[90] <= result_col4[89];
   result_col4[91] <= result_col4[90];
   result_col4[92] <= result_col4[91];
   result_col4[93] <= result_col4[92];
   result_col4[94] <= result_col4[93];
   result_col4[95] <= result_col4[94];
   result_col4[96] <= result_col4[95];
   result_col4[97] <= result_col4[96];
   result_col4[98] <= result_col4[97];
   result_col4[99] <= result_col4[98];
   result_col4[100] <= result_col4[99];
   result_col4[101] <= result_col4[100];
   result_col4[102] <= result_col4[101];
   result_col4[103] <= result_col4[102];
   result_col4[104] <= result_col4[103];
   result_col4[105] <= result_col4[104];
   result_col4[106] <= result_col4[105];
   result_col4[107] <= result_col4[106];
   result_col4[108] <= result_col4[107];
   result_col4[109] <= result_col4[108];
   result_col4[110] <= result_col4[109];
   result_col4[111] <= result_col4[110];
   result_col4[112] <= result_col4[111];
   result_col4[113] <= result_col4[112];
   result_col4[114] <= result_col4[113];
   result_col4[115] <= result_col4[114];
   result_col4[116] <= result_col4[115];
   result_col4[117] <= result_col4[116];
   result_col4[118] <= result_col4[117];
   result_col4[119] <= result_col4[118];
   result_col4[120] <= result_col4[119];
   result_col4[121] <= result_col4[120];
   result_col4[122] <= result_col4[121];
   result_col4[123] <= result_col4[122];
   result_col4[124] <= result_col4[123];
   result_col4[125] <= result_col4[124];
   result_col4[126] <= result_col4[125];
   result_col4[127] <= result_col4[126];
   result_col4[128] <= result_col4[127];
   result_col4[129] <= result_col4[128];
   result_col4[130] <= result_col4[129];
   result_col4[131] <= result_col4[130];
   result_col4[132] <= result_col4[131];
   result_col4[133] <= result_col4[132];
   result_col4[134] <= result_col4[133];
   result_col4[135] <= result_col4[134];
   result_col4[136] <= result_col4[135];
   result_col4[137] <= result_col4[136];
   result_col4[138] <= result_col4[137];
   result_col4[139] <= result_col4[138];
   result_col4[140] <= result_col4[139];
   result_col4[141] <= result_col4[140];
   result_col4[142] <= result_col4[141];
   result_col4[143] <= result_col4[142];
   result_col4[144] <= result_col4[143];
   result_col4[145] <= result_col4[144];
   result_col4[146] <= result_col4[145];
   result_col4[147] <= result_col4[146];
   result_col4[148] <= result_col4[147];
   result_col4[149] <= result_col4[148];
   result_col4[150] <= result_col4[149];
   result_col4[151] <= result_col4[150];
   result_col4[152] <= result_col4[151];
   result_col4[153] <= result_col4[152];
   result_col4[154] <= result_col4[153];
   result_col4[155] <= result_col4[154];
   result_col4[156] <= result_col4[155];
   result_col4[157] <= result_col4[156];
   result_col4[158] <= result_col4[157];
   result_col4[159] <= result_col4[158];
   result_col4[160] <= result_col4[159];
   result_col4[161] <= result_col4[160];
   result_col4[162] <= result_col4[161];

   result_col5[1] <= data_out_4_5;
   result_col5[2] <= result_col5[1];
   result_col5[3] <= result_col5[2];
   result_col5[4] <= result_col5[3];
   result_col5[5] <= result_col5[4];
   result_col5[6] <= result_col5[5];
   result_col5[7] <= result_col5[6];
   result_col5[8] <= result_col5[7];
   result_col5[9] <= result_col5[8];
   result_col5[10] <= result_col5[9];
   result_col5[11] <= result_col5[10];
   result_col5[12] <= result_col5[11];
   result_col5[13] <= result_col5[12];
   result_col5[14] <= result_col5[13];
   result_col5[15] <= result_col5[14];
   result_col5[16] <= result_col5[15];
   result_col5[17] <= result_col5[16];
   result_col5[18] <= result_col5[17];
   result_col5[19] <= result_col5[18];
   result_col5[20] <= result_col5[19];
   result_col5[21] <= result_col5[20];
   result_col5[22] <= result_col5[21];
   result_col5[23] <= result_col5[22];
   result_col5[24] <= result_col5[23];
   result_col5[25] <= result_col5[24];
   result_col5[26] <= result_col5[25];
   result_col5[27] <= result_col5[26];
   result_col5[28] <= result_col5[27];
   result_col5[29] <= result_col5[28];
   result_col5[30] <= result_col5[29];
   result_col5[31] <= result_col5[30];
   result_col5[32] <= result_col5[31];
   result_col5[33] <= result_col5[32];
   result_col5[34] <= result_col5[33];
   result_col5[35] <= result_col5[34];
   result_col5[36] <= result_col5[35];
   result_col5[37] <= result_col5[36];
   result_col5[38] <= result_col5[37];
   result_col5[39] <= result_col5[38];
   result_col5[40] <= result_col5[39];
   result_col5[41] <= result_col5[40];
   result_col5[42] <= result_col5[41];
   result_col5[43] <= result_col5[42];
   result_col5[44] <= result_col5[43];
   result_col5[45] <= result_col5[44];
   result_col5[46] <= result_col5[45];
   result_col5[47] <= result_col5[46];
   result_col5[48] <= result_col5[47];
   result_col5[49] <= result_col5[48];
   result_col5[50] <= result_col5[49];
   result_col5[51] <= result_col5[50];
   result_col5[52] <= result_col5[51];
   result_col5[53] <= result_col5[52];
   result_col5[54] <= result_col5[53];
   result_col5[55] <= result_col5[54];
   result_col5[56] <= result_col5[55];
   result_col5[57] <= result_col5[56];
   result_col5[58] <= result_col5[57];
   result_col5[59] <= result_col5[58];
   result_col5[60] <= result_col5[59];
   result_col5[61] <= result_col5[60];
   result_col5[62] <= result_col5[61];
   result_col5[63] <= result_col5[62];
   result_col5[64] <= result_col5[63];
   result_col5[65] <= result_col5[64];
   result_col5[66] <= result_col5[65];
   result_col5[67] <= result_col5[66];
   result_col5[68] <= result_col5[67];
   result_col5[69] <= result_col5[68];
   result_col5[70] <= result_col5[69];
   result_col5[71] <= result_col5[70];
   result_col5[72] <= result_col5[71];
   result_col5[73] <= result_col5[72];
   result_col5[74] <= result_col5[73];
   result_col5[75] <= result_col5[74];
   result_col5[76] <= result_col5[75];
   result_col5[77] <= result_col5[76];
   result_col5[78] <= result_col5[77];
   result_col5[79] <= result_col5[78];
   result_col5[80] <= result_col5[79];
   result_col5[81] <= result_col5[80];
   result_col5[82] <= result_col5[81];
   result_col5[83] <= result_col5[82];
   result_col5[84] <= result_col5[83];
   result_col5[85] <= result_col5[84];
   result_col5[86] <= result_col5[85];
   result_col5[87] <= result_col5[86];
   result_col5[88] <= result_col5[87];
   result_col5[89] <= result_col5[88];
   result_col5[90] <= result_col5[89];
   result_col5[91] <= result_col5[90];
   result_col5[92] <= result_col5[91];
   result_col5[93] <= result_col5[92];
   result_col5[94] <= result_col5[93];
   result_col5[95] <= result_col5[94];
   result_col5[96] <= result_col5[95];
   result_col5[97] <= result_col5[96];
   result_col5[98] <= result_col5[97];
   result_col5[99] <= result_col5[98];
   result_col5[100] <= result_col5[99];
   result_col5[101] <= result_col5[100];
   result_col5[102] <= result_col5[101];
   result_col5[103] <= result_col5[102];
   result_col5[104] <= result_col5[103];
   result_col5[105] <= result_col5[104];
   result_col5[106] <= result_col5[105];
   result_col5[107] <= result_col5[106];
   result_col5[108] <= result_col5[107];
   result_col5[109] <= result_col5[108];
   result_col5[110] <= result_col5[109];
   result_col5[111] <= result_col5[110];
   result_col5[112] <= result_col5[111];
   result_col5[113] <= result_col5[112];
   result_col5[114] <= result_col5[113];
   result_col5[115] <= result_col5[114];
   result_col5[116] <= result_col5[115];
   result_col5[117] <= result_col5[116];
   result_col5[118] <= result_col5[117];
   result_col5[119] <= result_col5[118];
   result_col5[120] <= result_col5[119];
   result_col5[121] <= result_col5[120];
   result_col5[122] <= result_col5[121];
   result_col5[123] <= result_col5[122];
   result_col5[124] <= result_col5[123];
   result_col5[125] <= result_col5[124];
   result_col5[126] <= result_col5[125];
   result_col5[127] <= result_col5[126];
   result_col5[128] <= result_col5[127];
   result_col5[129] <= result_col5[128];
   result_col5[130] <= result_col5[129];
   result_col5[131] <= result_col5[130];
   result_col5[132] <= result_col5[131];
   result_col5[133] <= result_col5[132];
   result_col5[134] <= result_col5[133];
   result_col5[135] <= result_col5[134];
   result_col5[136] <= result_col5[135];
   result_col5[137] <= result_col5[136];
   result_col5[138] <= result_col5[137];
   result_col5[139] <= result_col5[138];
   result_col5[140] <= result_col5[139];
   result_col5[141] <= result_col5[140];
   result_col5[142] <= result_col5[141];
   result_col5[143] <= result_col5[142];
   result_col5[144] <= result_col5[143];
   result_col5[145] <= result_col5[144];
   result_col5[146] <= result_col5[145];
   result_col5[147] <= result_col5[146];
   result_col5[148] <= result_col5[147];
   result_col5[149] <= result_col5[148];
   result_col5[150] <= result_col5[149];
   result_col5[151] <= result_col5[150];
   result_col5[152] <= result_col5[151];
   result_col5[153] <= result_col5[152];
   result_col5[154] <= result_col5[153];
   result_col5[155] <= result_col5[154];
   result_col5[156] <= result_col5[155];
   result_col5[157] <= result_col5[156];
   result_col5[158] <= result_col5[157];
   result_col5[159] <= result_col5[158];
   result_col5[160] <= result_col5[159];
   result_col5[161] <= result_col5[160];

   result_col6[1] <= data_out_4_6;
   result_col6[2] <= result_col6[1];
   result_col6[3] <= result_col6[2];
   result_col6[4] <= result_col6[3];
   result_col6[5] <= result_col6[4];
   result_col6[6] <= result_col6[5];
   result_col6[7] <= result_col6[6];
   result_col6[8] <= result_col6[7];
   result_col6[9] <= result_col6[8];
   result_col6[10] <= result_col6[9];
   result_col6[11] <= result_col6[10];
   result_col6[12] <= result_col6[11];
   result_col6[13] <= result_col6[12];
   result_col6[14] <= result_col6[13];
   result_col6[15] <= result_col6[14];
   result_col6[16] <= result_col6[15];
   result_col6[17] <= result_col6[16];
   result_col6[18] <= result_col6[17];
   result_col6[19] <= result_col6[18];
   result_col6[20] <= result_col6[19];
   result_col6[21] <= result_col6[20];
   result_col6[22] <= result_col6[21];
   result_col6[23] <= result_col6[22];
   result_col6[24] <= result_col6[23];
   result_col6[25] <= result_col6[24];
   result_col6[26] <= result_col6[25];
   result_col6[27] <= result_col6[26];
   result_col6[28] <= result_col6[27];
   result_col6[29] <= result_col6[28];
   result_col6[30] <= result_col6[29];
   result_col6[31] <= result_col6[30];
   result_col6[32] <= result_col6[31];
   result_col6[33] <= result_col6[32];
   result_col6[34] <= result_col6[33];
   result_col6[35] <= result_col6[34];
   result_col6[36] <= result_col6[35];
   result_col6[37] <= result_col6[36];
   result_col6[38] <= result_col6[37];
   result_col6[39] <= result_col6[38];
   result_col6[40] <= result_col6[39];
   result_col6[41] <= result_col6[40];
   result_col6[42] <= result_col6[41];
   result_col6[43] <= result_col6[42];
   result_col6[44] <= result_col6[43];
   result_col6[45] <= result_col6[44];
   result_col6[46] <= result_col6[45];
   result_col6[47] <= result_col6[46];
   result_col6[48] <= result_col6[47];
   result_col6[49] <= result_col6[48];
   result_col6[50] <= result_col6[49];
   result_col6[51] <= result_col6[50];
   result_col6[52] <= result_col6[51];
   result_col6[53] <= result_col6[52];
   result_col6[54] <= result_col6[53];
   result_col6[55] <= result_col6[54];
   result_col6[56] <= result_col6[55];
   result_col6[57] <= result_col6[56];
   result_col6[58] <= result_col6[57];
   result_col6[59] <= result_col6[58];
   result_col6[60] <= result_col6[59];
   result_col6[61] <= result_col6[60];
   result_col6[62] <= result_col6[61];
   result_col6[63] <= result_col6[62];
   result_col6[64] <= result_col6[63];
   result_col6[65] <= result_col6[64];
   result_col6[66] <= result_col6[65];
   result_col6[67] <= result_col6[66];
   result_col6[68] <= result_col6[67];
   result_col6[69] <= result_col6[68];
   result_col6[70] <= result_col6[69];
   result_col6[71] <= result_col6[70];
   result_col6[72] <= result_col6[71];
   result_col6[73] <= result_col6[72];
   result_col6[74] <= result_col6[73];
   result_col6[75] <= result_col6[74];
   result_col6[76] <= result_col6[75];
   result_col6[77] <= result_col6[76];
   result_col6[78] <= result_col6[77];
   result_col6[79] <= result_col6[78];
   result_col6[80] <= result_col6[79];
   result_col6[81] <= result_col6[80];
   result_col6[82] <= result_col6[81];
   result_col6[83] <= result_col6[82];
   result_col6[84] <= result_col6[83];
   result_col6[85] <= result_col6[84];
   result_col6[86] <= result_col6[85];
   result_col6[87] <= result_col6[86];
   result_col6[88] <= result_col6[87];
   result_col6[89] <= result_col6[88];
   result_col6[90] <= result_col6[89];
   result_col6[91] <= result_col6[90];
   result_col6[92] <= result_col6[91];
   result_col6[93] <= result_col6[92];
   result_col6[94] <= result_col6[93];
   result_col6[95] <= result_col6[94];
   result_col6[96] <= result_col6[95];
   result_col6[97] <= result_col6[96];
   result_col6[98] <= result_col6[97];
   result_col6[99] <= result_col6[98];
   result_col6[100] <= result_col6[99];
   result_col6[101] <= result_col6[100];
   result_col6[102] <= result_col6[101];
   result_col6[103] <= result_col6[102];
   result_col6[104] <= result_col6[103];
   result_col6[105] <= result_col6[104];
   result_col6[106] <= result_col6[105];
   result_col6[107] <= result_col6[106];
   result_col6[108] <= result_col6[107];
   result_col6[109] <= result_col6[108];
   result_col6[110] <= result_col6[109];
   result_col6[111] <= result_col6[110];
   result_col6[112] <= result_col6[111];
   result_col6[113] <= result_col6[112];
   result_col6[114] <= result_col6[113];
   result_col6[115] <= result_col6[114];
   result_col6[116] <= result_col6[115];
   result_col6[117] <= result_col6[116];
   result_col6[118] <= result_col6[117];
   result_col6[119] <= result_col6[118];
   result_col6[120] <= result_col6[119];
   result_col6[121] <= result_col6[120];
   result_col6[122] <= result_col6[121];
   result_col6[123] <= result_col6[122];
   result_col6[124] <= result_col6[123];
   result_col6[125] <= result_col6[124];
   result_col6[126] <= result_col6[125];
   result_col6[127] <= result_col6[126];
   result_col6[128] <= result_col6[127];
   result_col6[129] <= result_col6[128];
   result_col6[130] <= result_col6[129];
   result_col6[131] <= result_col6[130];
   result_col6[132] <= result_col6[131];
   result_col6[133] <= result_col6[132];
   result_col6[134] <= result_col6[133];
   result_col6[135] <= result_col6[134];
   result_col6[136] <= result_col6[135];
   result_col6[137] <= result_col6[136];
   result_col6[138] <= result_col6[137];
   result_col6[139] <= result_col6[138];
   result_col6[140] <= result_col6[139];
   result_col6[141] <= result_col6[140];
   result_col6[142] <= result_col6[141];
   result_col6[143] <= result_col6[142];
   result_col6[144] <= result_col6[143];
   result_col6[145] <= result_col6[144];
   result_col6[146] <= result_col6[145];
   result_col6[147] <= result_col6[146];
   result_col6[148] <= result_col6[147];
   result_col6[149] <= result_col6[148];
   result_col6[150] <= result_col6[149];
   result_col6[151] <= result_col6[150];
   result_col6[152] <= result_col6[151];
   result_col6[153] <= result_col6[152];
   result_col6[154] <= result_col6[153];
   result_col6[155] <= result_col6[154];
   result_col6[156] <= result_col6[155];
   result_col6[157] <= result_col6[156];
   result_col6[158] <= result_col6[157];
   result_col6[159] <= result_col6[158];
   result_col6[160] <= result_col6[159];

   result_col7[1] <= data_out_4_7;
   result_col7[2] <= result_col7[1];
   result_col7[3] <= result_col7[2];
   result_col7[4] <= result_col7[3];
   result_col7[5] <= result_col7[4];
   result_col7[6] <= result_col7[5];
   result_col7[7] <= result_col7[6];
   result_col7[8] <= result_col7[7];
   result_col7[9] <= result_col7[8];
   result_col7[10] <= result_col7[9];
   result_col7[11] <= result_col7[10];
   result_col7[12] <= result_col7[11];
   result_col7[13] <= result_col7[12];
   result_col7[14] <= result_col7[13];
   result_col7[15] <= result_col7[14];
   result_col7[16] <= result_col7[15];
   result_col7[17] <= result_col7[16];
   result_col7[18] <= result_col7[17];
   result_col7[19] <= result_col7[18];
   result_col7[20] <= result_col7[19];
   result_col7[21] <= result_col7[20];
   result_col7[22] <= result_col7[21];
   result_col7[23] <= result_col7[22];
   result_col7[24] <= result_col7[23];
   result_col7[25] <= result_col7[24];
   result_col7[26] <= result_col7[25];
   result_col7[27] <= result_col7[26];
   result_col7[28] <= result_col7[27];
   result_col7[29] <= result_col7[28];
   result_col7[30] <= result_col7[29];
   result_col7[31] <= result_col7[30];
   result_col7[32] <= result_col7[31];
   result_col7[33] <= result_col7[32];
   result_col7[34] <= result_col7[33];
   result_col7[35] <= result_col7[34];
   result_col7[36] <= result_col7[35];
   result_col7[37] <= result_col7[36];
   result_col7[38] <= result_col7[37];
   result_col7[39] <= result_col7[38];
   result_col7[40] <= result_col7[39];
   result_col7[41] <= result_col7[40];
   result_col7[42] <= result_col7[41];
   result_col7[43] <= result_col7[42];
   result_col7[44] <= result_col7[43];
   result_col7[45] <= result_col7[44];
   result_col7[46] <= result_col7[45];
   result_col7[47] <= result_col7[46];
   result_col7[48] <= result_col7[47];
   result_col7[49] <= result_col7[48];
   result_col7[50] <= result_col7[49];
   result_col7[51] <= result_col7[50];
   result_col7[52] <= result_col7[51];
   result_col7[53] <= result_col7[52];
   result_col7[54] <= result_col7[53];
   result_col7[55] <= result_col7[54];
   result_col7[56] <= result_col7[55];
   result_col7[57] <= result_col7[56];
   result_col7[58] <= result_col7[57];
   result_col7[59] <= result_col7[58];
   result_col7[60] <= result_col7[59];
   result_col7[61] <= result_col7[60];
   result_col7[62] <= result_col7[61];
   result_col7[63] <= result_col7[62];
   result_col7[64] <= result_col7[63];
   result_col7[65] <= result_col7[64];
   result_col7[66] <= result_col7[65];
   result_col7[67] <= result_col7[66];
   result_col7[68] <= result_col7[67];
   result_col7[69] <= result_col7[68];
   result_col7[70] <= result_col7[69];
   result_col7[71] <= result_col7[70];
   result_col7[72] <= result_col7[71];
   result_col7[73] <= result_col7[72];
   result_col7[74] <= result_col7[73];
   result_col7[75] <= result_col7[74];
   result_col7[76] <= result_col7[75];
   result_col7[77] <= result_col7[76];
   result_col7[78] <= result_col7[77];
   result_col7[79] <= result_col7[78];
   result_col7[80] <= result_col7[79];
   result_col7[81] <= result_col7[80];
   result_col7[82] <= result_col7[81];
   result_col7[83] <= result_col7[82];
   result_col7[84] <= result_col7[83];
   result_col7[85] <= result_col7[84];
   result_col7[86] <= result_col7[85];
   result_col7[87] <= result_col7[86];
   result_col7[88] <= result_col7[87];
   result_col7[89] <= result_col7[88];
   result_col7[90] <= result_col7[89];
   result_col7[91] <= result_col7[90];
   result_col7[92] <= result_col7[91];
   result_col7[93] <= result_col7[92];
   result_col7[94] <= result_col7[93];
   result_col7[95] <= result_col7[94];
   result_col7[96] <= result_col7[95];
   result_col7[97] <= result_col7[96];
   result_col7[98] <= result_col7[97];
   result_col7[99] <= result_col7[98];
   result_col7[100] <= result_col7[99];
   result_col7[101] <= result_col7[100];
   result_col7[102] <= result_col7[101];
   result_col7[103] <= result_col7[102];
   result_col7[104] <= result_col7[103];
   result_col7[105] <= result_col7[104];
   result_col7[106] <= result_col7[105];
   result_col7[107] <= result_col7[106];
   result_col7[108] <= result_col7[107];
   result_col7[109] <= result_col7[108];
   result_col7[110] <= result_col7[109];
   result_col7[111] <= result_col7[110];
   result_col7[112] <= result_col7[111];
   result_col7[113] <= result_col7[112];
   result_col7[114] <= result_col7[113];
   result_col7[115] <= result_col7[114];
   result_col7[116] <= result_col7[115];
   result_col7[117] <= result_col7[116];
   result_col7[118] <= result_col7[117];
   result_col7[119] <= result_col7[118];
   result_col7[120] <= result_col7[119];
   result_col7[121] <= result_col7[120];
   result_col7[122] <= result_col7[121];
   result_col7[123] <= result_col7[122];
   result_col7[124] <= result_col7[123];
   result_col7[125] <= result_col7[124];
   result_col7[126] <= result_col7[125];
   result_col7[127] <= result_col7[126];
   result_col7[128] <= result_col7[127];
   result_col7[129] <= result_col7[128];
   result_col7[130] <= result_col7[129];
   result_col7[131] <= result_col7[130];
   result_col7[132] <= result_col7[131];
   result_col7[133] <= result_col7[132];
   result_col7[134] <= result_col7[133];
   result_col7[135] <= result_col7[134];
   result_col7[136] <= result_col7[135];
   result_col7[137] <= result_col7[136];
   result_col7[138] <= result_col7[137];
   result_col7[139] <= result_col7[138];
   result_col7[140] <= result_col7[139];
   result_col7[141] <= result_col7[140];
   result_col7[142] <= result_col7[141];
   result_col7[143] <= result_col7[142];
   result_col7[144] <= result_col7[143];
   result_col7[145] <= result_col7[144];
   result_col7[146] <= result_col7[145];
   result_col7[147] <= result_col7[146];
   result_col7[148] <= result_col7[147];
   result_col7[149] <= result_col7[148];
   result_col7[150] <= result_col7[149];
   result_col7[151] <= result_col7[150];
   result_col7[152] <= result_col7[151];
   result_col7[153] <= result_col7[152];
   result_col7[154] <= result_col7[153];
   result_col7[155] <= result_col7[154];
   result_col7[156] <= result_col7[155];
   result_col7[157] <= result_col7[156];
   result_col7[158] <= result_col7[157];
   result_col7[159] <= result_col7[158];

   result_col8[1] <= data_out_4_8;
   result_col8[2] <= result_col8[1];
   result_col8[3] <= result_col8[2];
   result_col8[4] <= result_col8[3];
   result_col8[5] <= result_col8[4];
   result_col8[6] <= result_col8[5];
   result_col8[7] <= result_col8[6];
   result_col8[8] <= result_col8[7];
   result_col8[9] <= result_col8[8];
   result_col8[10] <= result_col8[9];
   result_col8[11] <= result_col8[10];
   result_col8[12] <= result_col8[11];
   result_col8[13] <= result_col8[12];
   result_col8[14] <= result_col8[13];
   result_col8[15] <= result_col8[14];
   result_col8[16] <= result_col8[15];
   result_col8[17] <= result_col8[16];
   result_col8[18] <= result_col8[17];
   result_col8[19] <= result_col8[18];
   result_col8[20] <= result_col8[19];
   result_col8[21] <= result_col8[20];
   result_col8[22] <= result_col8[21];
   result_col8[23] <= result_col8[22];
   result_col8[24] <= result_col8[23];
   result_col8[25] <= result_col8[24];
   result_col8[26] <= result_col8[25];
   result_col8[27] <= result_col8[26];
   result_col8[28] <= result_col8[27];
   result_col8[29] <= result_col8[28];
   result_col8[30] <= result_col8[29];
   result_col8[31] <= result_col8[30];
   result_col8[32] <= result_col8[31];
   result_col8[33] <= result_col8[32];
   result_col8[34] <= result_col8[33];
   result_col8[35] <= result_col8[34];
   result_col8[36] <= result_col8[35];
   result_col8[37] <= result_col8[36];
   result_col8[38] <= result_col8[37];
   result_col8[39] <= result_col8[38];
   result_col8[40] <= result_col8[39];
   result_col8[41] <= result_col8[40];
   result_col8[42] <= result_col8[41];
   result_col8[43] <= result_col8[42];
   result_col8[44] <= result_col8[43];
   result_col8[45] <= result_col8[44];
   result_col8[46] <= result_col8[45];
   result_col8[47] <= result_col8[46];
   result_col8[48] <= result_col8[47];
   result_col8[49] <= result_col8[48];
   result_col8[50] <= result_col8[49];
   result_col8[51] <= result_col8[50];
   result_col8[52] <= result_col8[51];
   result_col8[53] <= result_col8[52];
   result_col8[54] <= result_col8[53];
   result_col8[55] <= result_col8[54];
   result_col8[56] <= result_col8[55];
   result_col8[57] <= result_col8[56];
   result_col8[58] <= result_col8[57];
   result_col8[59] <= result_col8[58];
   result_col8[60] <= result_col8[59];
   result_col8[61] <= result_col8[60];
   result_col8[62] <= result_col8[61];
   result_col8[63] <= result_col8[62];
   result_col8[64] <= result_col8[63];
   result_col8[65] <= result_col8[64];
   result_col8[66] <= result_col8[65];
   result_col8[67] <= result_col8[66];
   result_col8[68] <= result_col8[67];
   result_col8[69] <= result_col8[68];
   result_col8[70] <= result_col8[69];
   result_col8[71] <= result_col8[70];
   result_col8[72] <= result_col8[71];
   result_col8[73] <= result_col8[72];
   result_col8[74] <= result_col8[73];
   result_col8[75] <= result_col8[74];
   result_col8[76] <= result_col8[75];
   result_col8[77] <= result_col8[76];
   result_col8[78] <= result_col8[77];
   result_col8[79] <= result_col8[78];
   result_col8[80] <= result_col8[79];
   result_col8[81] <= result_col8[80];
   result_col8[82] <= result_col8[81];
   result_col8[83] <= result_col8[82];
   result_col8[84] <= result_col8[83];
   result_col8[85] <= result_col8[84];
   result_col8[86] <= result_col8[85];
   result_col8[87] <= result_col8[86];
   result_col8[88] <= result_col8[87];
   result_col8[89] <= result_col8[88];
   result_col8[90] <= result_col8[89];
   result_col8[91] <= result_col8[90];
   result_col8[92] <= result_col8[91];
   result_col8[93] <= result_col8[92];
   result_col8[94] <= result_col8[93];
   result_col8[95] <= result_col8[94];
   result_col8[96] <= result_col8[95];
   result_col8[97] <= result_col8[96];
   result_col8[98] <= result_col8[97];
   result_col8[99] <= result_col8[98];
   result_col8[100] <= result_col8[99];
   result_col8[101] <= result_col8[100];
   result_col8[102] <= result_col8[101];
   result_col8[103] <= result_col8[102];
   result_col8[104] <= result_col8[103];
   result_col8[105] <= result_col8[104];
   result_col8[106] <= result_col8[105];
   result_col8[107] <= result_col8[106];
   result_col8[108] <= result_col8[107];
   result_col8[109] <= result_col8[108];
   result_col8[110] <= result_col8[109];
   result_col8[111] <= result_col8[110];
   result_col8[112] <= result_col8[111];
   result_col8[113] <= result_col8[112];
   result_col8[114] <= result_col8[113];
   result_col8[115] <= result_col8[114];
   result_col8[116] <= result_col8[115];
   result_col8[117] <= result_col8[116];
   result_col8[118] <= result_col8[117];
   result_col8[119] <= result_col8[118];
   result_col8[120] <= result_col8[119];
   result_col8[121] <= result_col8[120];
   result_col8[122] <= result_col8[121];
   result_col8[123] <= result_col8[122];
   result_col8[124] <= result_col8[123];
   result_col8[125] <= result_col8[124];
   result_col8[126] <= result_col8[125];
   result_col8[127] <= result_col8[126];
   result_col8[128] <= result_col8[127];
   result_col8[129] <= result_col8[128];
   result_col8[130] <= result_col8[129];
   result_col8[131] <= result_col8[130];
   result_col8[132] <= result_col8[131];
   result_col8[133] <= result_col8[132];
   result_col8[134] <= result_col8[133];
   result_col8[135] <= result_col8[134];
   result_col8[136] <= result_col8[135];
   result_col8[137] <= result_col8[136];
   result_col8[138] <= result_col8[137];
   result_col8[139] <= result_col8[138];
   result_col8[140] <= result_col8[139];
   result_col8[141] <= result_col8[140];
   result_col8[142] <= result_col8[141];
   result_col8[143] <= result_col8[142];
   result_col8[144] <= result_col8[143];
   result_col8[145] <= result_col8[144];
   result_col8[146] <= result_col8[145];
   result_col8[147] <= result_col8[146];
   result_col8[148] <= result_col8[147];
   result_col8[149] <= result_col8[148];
   result_col8[150] <= result_col8[149];
   result_col8[151] <= result_col8[150];
   result_col8[152] <= result_col8[151];
   result_col8[153] <= result_col8[152];
   result_col8[154] <= result_col8[153];
   result_col8[155] <= result_col8[154];
   result_col8[156] <= result_col8[155];
   result_col8[157] <= result_col8[156];
   result_col8[158] <= result_col8[157];

   result_col9[1] <= data_out_4_9;
   result_col9[2] <= result_col9[1];
   result_col9[3] <= result_col9[2];
   result_col9[4] <= result_col9[3];
   result_col9[5] <= result_col9[4];
   result_col9[6] <= result_col9[5];
   result_col9[7] <= result_col9[6];
   result_col9[8] <= result_col9[7];
   result_col9[9] <= result_col9[8];
   result_col9[10] <= result_col9[9];
   result_col9[11] <= result_col9[10];
   result_col9[12] <= result_col9[11];
   result_col9[13] <= result_col9[12];
   result_col9[14] <= result_col9[13];
   result_col9[15] <= result_col9[14];
   result_col9[16] <= result_col9[15];
   result_col9[17] <= result_col9[16];
   result_col9[18] <= result_col9[17];
   result_col9[19] <= result_col9[18];
   result_col9[20] <= result_col9[19];
   result_col9[21] <= result_col9[20];
   result_col9[22] <= result_col9[21];
   result_col9[23] <= result_col9[22];
   result_col9[24] <= result_col9[23];
   result_col9[25] <= result_col9[24];
   result_col9[26] <= result_col9[25];
   result_col9[27] <= result_col9[26];
   result_col9[28] <= result_col9[27];
   result_col9[29] <= result_col9[28];
   result_col9[30] <= result_col9[29];
   result_col9[31] <= result_col9[30];
   result_col9[32] <= result_col9[31];
   result_col9[33] <= result_col9[32];
   result_col9[34] <= result_col9[33];
   result_col9[35] <= result_col9[34];
   result_col9[36] <= result_col9[35];
   result_col9[37] <= result_col9[36];
   result_col9[38] <= result_col9[37];
   result_col9[39] <= result_col9[38];
   result_col9[40] <= result_col9[39];
   result_col9[41] <= result_col9[40];
   result_col9[42] <= result_col9[41];
   result_col9[43] <= result_col9[42];
   result_col9[44] <= result_col9[43];
   result_col9[45] <= result_col9[44];
   result_col9[46] <= result_col9[45];
   result_col9[47] <= result_col9[46];
   result_col9[48] <= result_col9[47];
   result_col9[49] <= result_col9[48];
   result_col9[50] <= result_col9[49];
   result_col9[51] <= result_col9[50];
   result_col9[52] <= result_col9[51];
   result_col9[53] <= result_col9[52];
   result_col9[54] <= result_col9[53];
   result_col9[55] <= result_col9[54];
   result_col9[56] <= result_col9[55];
   result_col9[57] <= result_col9[56];
   result_col9[58] <= result_col9[57];
   result_col9[59] <= result_col9[58];
   result_col9[60] <= result_col9[59];
   result_col9[61] <= result_col9[60];
   result_col9[62] <= result_col9[61];
   result_col9[63] <= result_col9[62];
   result_col9[64] <= result_col9[63];
   result_col9[65] <= result_col9[64];
   result_col9[66] <= result_col9[65];
   result_col9[67] <= result_col9[66];
   result_col9[68] <= result_col9[67];
   result_col9[69] <= result_col9[68];
   result_col9[70] <= result_col9[69];
   result_col9[71] <= result_col9[70];
   result_col9[72] <= result_col9[71];
   result_col9[73] <= result_col9[72];
   result_col9[74] <= result_col9[73];
   result_col9[75] <= result_col9[74];
   result_col9[76] <= result_col9[75];
   result_col9[77] <= result_col9[76];
   result_col9[78] <= result_col9[77];
   result_col9[79] <= result_col9[78];
   result_col9[80] <= result_col9[79];
   result_col9[81] <= result_col9[80];
   result_col9[82] <= result_col9[81];
   result_col9[83] <= result_col9[82];
   result_col9[84] <= result_col9[83];
   result_col9[85] <= result_col9[84];
   result_col9[86] <= result_col9[85];
   result_col9[87] <= result_col9[86];
   result_col9[88] <= result_col9[87];
   result_col9[89] <= result_col9[88];
   result_col9[90] <= result_col9[89];
   result_col9[91] <= result_col9[90];
   result_col9[92] <= result_col9[91];
   result_col9[93] <= result_col9[92];
   result_col9[94] <= result_col9[93];
   result_col9[95] <= result_col9[94];
   result_col9[96] <= result_col9[95];
   result_col9[97] <= result_col9[96];
   result_col9[98] <= result_col9[97];
   result_col9[99] <= result_col9[98];
   result_col9[100] <= result_col9[99];
   result_col9[101] <= result_col9[100];
   result_col9[102] <= result_col9[101];
   result_col9[103] <= result_col9[102];
   result_col9[104] <= result_col9[103];
   result_col9[105] <= result_col9[104];
   result_col9[106] <= result_col9[105];
   result_col9[107] <= result_col9[106];
   result_col9[108] <= result_col9[107];
   result_col9[109] <= result_col9[108];
   result_col9[110] <= result_col9[109];
   result_col9[111] <= result_col9[110];
   result_col9[112] <= result_col9[111];
   result_col9[113] <= result_col9[112];
   result_col9[114] <= result_col9[113];
   result_col9[115] <= result_col9[114];
   result_col9[116] <= result_col9[115];
   result_col9[117] <= result_col9[116];
   result_col9[118] <= result_col9[117];
   result_col9[119] <= result_col9[118];
   result_col9[120] <= result_col9[119];
   result_col9[121] <= result_col9[120];
   result_col9[122] <= result_col9[121];
   result_col9[123] <= result_col9[122];
   result_col9[124] <= result_col9[123];
   result_col9[125] <= result_col9[124];
   result_col9[126] <= result_col9[125];
   result_col9[127] <= result_col9[126];
   result_col9[128] <= result_col9[127];
   result_col9[129] <= result_col9[128];
   result_col9[130] <= result_col9[129];
   result_col9[131] <= result_col9[130];
   result_col9[132] <= result_col9[131];
   result_col9[133] <= result_col9[132];
   result_col9[134] <= result_col9[133];
   result_col9[135] <= result_col9[134];
   result_col9[136] <= result_col9[135];
   result_col9[137] <= result_col9[136];
   result_col9[138] <= result_col9[137];
   result_col9[139] <= result_col9[138];
   result_col9[140] <= result_col9[139];
   result_col9[141] <= result_col9[140];
   result_col9[142] <= result_col9[141];
   result_col9[143] <= result_col9[142];
   result_col9[144] <= result_col9[143];
   result_col9[145] <= result_col9[144];
   result_col9[146] <= result_col9[145];
   result_col9[147] <= result_col9[146];
   result_col9[148] <= result_col9[147];
   result_col9[149] <= result_col9[148];
   result_col9[150] <= result_col9[149];
   result_col9[151] <= result_col9[150];
   result_col9[152] <= result_col9[151];
   result_col9[153] <= result_col9[152];
   result_col9[154] <= result_col9[153];
   result_col9[155] <= result_col9[154];
   result_col9[156] <= result_col9[155];
   result_col9[157] <= result_col9[156];

   result_col10[1] <= data_out_4_10;
   result_col10[2] <= result_col10[1];
   result_col10[3] <= result_col10[2];
   result_col10[4] <= result_col10[3];
   result_col10[5] <= result_col10[4];
   result_col10[6] <= result_col10[5];
   result_col10[7] <= result_col10[6];
   result_col10[8] <= result_col10[7];
   result_col10[9] <= result_col10[8];
   result_col10[10] <= result_col10[9];
   result_col10[11] <= result_col10[10];
   result_col10[12] <= result_col10[11];
   result_col10[13] <= result_col10[12];
   result_col10[14] <= result_col10[13];
   result_col10[15] <= result_col10[14];
   result_col10[16] <= result_col10[15];
   result_col10[17] <= result_col10[16];
   result_col10[18] <= result_col10[17];
   result_col10[19] <= result_col10[18];
   result_col10[20] <= result_col10[19];
   result_col10[21] <= result_col10[20];
   result_col10[22] <= result_col10[21];
   result_col10[23] <= result_col10[22];
   result_col10[24] <= result_col10[23];
   result_col10[25] <= result_col10[24];
   result_col10[26] <= result_col10[25];
   result_col10[27] <= result_col10[26];
   result_col10[28] <= result_col10[27];
   result_col10[29] <= result_col10[28];
   result_col10[30] <= result_col10[29];
   result_col10[31] <= result_col10[30];
   result_col10[32] <= result_col10[31];
   result_col10[33] <= result_col10[32];
   result_col10[34] <= result_col10[33];
   result_col10[35] <= result_col10[34];
   result_col10[36] <= result_col10[35];
   result_col10[37] <= result_col10[36];
   result_col10[38] <= result_col10[37];
   result_col10[39] <= result_col10[38];
   result_col10[40] <= result_col10[39];
   result_col10[41] <= result_col10[40];
   result_col10[42] <= result_col10[41];
   result_col10[43] <= result_col10[42];
   result_col10[44] <= result_col10[43];
   result_col10[45] <= result_col10[44];
   result_col10[46] <= result_col10[45];
   result_col10[47] <= result_col10[46];
   result_col10[48] <= result_col10[47];
   result_col10[49] <= result_col10[48];
   result_col10[50] <= result_col10[49];
   result_col10[51] <= result_col10[50];
   result_col10[52] <= result_col10[51];
   result_col10[53] <= result_col10[52];
   result_col10[54] <= result_col10[53];
   result_col10[55] <= result_col10[54];
   result_col10[56] <= result_col10[55];
   result_col10[57] <= result_col10[56];
   result_col10[58] <= result_col10[57];
   result_col10[59] <= result_col10[58];
   result_col10[60] <= result_col10[59];
   result_col10[61] <= result_col10[60];
   result_col10[62] <= result_col10[61];
   result_col10[63] <= result_col10[62];
   result_col10[64] <= result_col10[63];
   result_col10[65] <= result_col10[64];
   result_col10[66] <= result_col10[65];
   result_col10[67] <= result_col10[66];
   result_col10[68] <= result_col10[67];
   result_col10[69] <= result_col10[68];
   result_col10[70] <= result_col10[69];
   result_col10[71] <= result_col10[70];
   result_col10[72] <= result_col10[71];
   result_col10[73] <= result_col10[72];
   result_col10[74] <= result_col10[73];
   result_col10[75] <= result_col10[74];
   result_col10[76] <= result_col10[75];
   result_col10[77] <= result_col10[76];
   result_col10[78] <= result_col10[77];
   result_col10[79] <= result_col10[78];
   result_col10[80] <= result_col10[79];
   result_col10[81] <= result_col10[80];
   result_col10[82] <= result_col10[81];
   result_col10[83] <= result_col10[82];
   result_col10[84] <= result_col10[83];
   result_col10[85] <= result_col10[84];
   result_col10[86] <= result_col10[85];
   result_col10[87] <= result_col10[86];
   result_col10[88] <= result_col10[87];
   result_col10[89] <= result_col10[88];
   result_col10[90] <= result_col10[89];
   result_col10[91] <= result_col10[90];
   result_col10[92] <= result_col10[91];
   result_col10[93] <= result_col10[92];
   result_col10[94] <= result_col10[93];
   result_col10[95] <= result_col10[94];
   result_col10[96] <= result_col10[95];
   result_col10[97] <= result_col10[96];
   result_col10[98] <= result_col10[97];
   result_col10[99] <= result_col10[98];
   result_col10[100] <= result_col10[99];
   result_col10[101] <= result_col10[100];
   result_col10[102] <= result_col10[101];
   result_col10[103] <= result_col10[102];
   result_col10[104] <= result_col10[103];
   result_col10[105] <= result_col10[104];
   result_col10[106] <= result_col10[105];
   result_col10[107] <= result_col10[106];
   result_col10[108] <= result_col10[107];
   result_col10[109] <= result_col10[108];
   result_col10[110] <= result_col10[109];
   result_col10[111] <= result_col10[110];
   result_col10[112] <= result_col10[111];
   result_col10[113] <= result_col10[112];
   result_col10[114] <= result_col10[113];
   result_col10[115] <= result_col10[114];
   result_col10[116] <= result_col10[115];
   result_col10[117] <= result_col10[116];
   result_col10[118] <= result_col10[117];
   result_col10[119] <= result_col10[118];
   result_col10[120] <= result_col10[119];
   result_col10[121] <= result_col10[120];
   result_col10[122] <= result_col10[121];
   result_col10[123] <= result_col10[122];
   result_col10[124] <= result_col10[123];
   result_col10[125] <= result_col10[124];
   result_col10[126] <= result_col10[125];
   result_col10[127] <= result_col10[126];
   result_col10[128] <= result_col10[127];
   result_col10[129] <= result_col10[128];
   result_col10[130] <= result_col10[129];
   result_col10[131] <= result_col10[130];
   result_col10[132] <= result_col10[131];
   result_col10[133] <= result_col10[132];
   result_col10[134] <= result_col10[133];
   result_col10[135] <= result_col10[134];
   result_col10[136] <= result_col10[135];
   result_col10[137] <= result_col10[136];
   result_col10[138] <= result_col10[137];
   result_col10[139] <= result_col10[138];
   result_col10[140] <= result_col10[139];
   result_col10[141] <= result_col10[140];
   result_col10[142] <= result_col10[141];
   result_col10[143] <= result_col10[142];
   result_col10[144] <= result_col10[143];
   result_col10[145] <= result_col10[144];
   result_col10[146] <= result_col10[145];
   result_col10[147] <= result_col10[146];
   result_col10[148] <= result_col10[147];
   result_col10[149] <= result_col10[148];
   result_col10[150] <= result_col10[149];
   result_col10[151] <= result_col10[150];
   result_col10[152] <= result_col10[151];
   result_col10[153] <= result_col10[152];
   result_col10[154] <= result_col10[153];
   result_col10[155] <= result_col10[154];
   result_col10[156] <= result_col10[155];

   result_col11[1] <= data_out_4_11;
   result_col11[2] <= result_col11[1];
   result_col11[3] <= result_col11[2];
   result_col11[4] <= result_col11[3];
   result_col11[5] <= result_col11[4];
   result_col11[6] <= result_col11[5];
   result_col11[7] <= result_col11[6];
   result_col11[8] <= result_col11[7];
   result_col11[9] <= result_col11[8];
   result_col11[10] <= result_col11[9];
   result_col11[11] <= result_col11[10];
   result_col11[12] <= result_col11[11];
   result_col11[13] <= result_col11[12];
   result_col11[14] <= result_col11[13];
   result_col11[15] <= result_col11[14];
   result_col11[16] <= result_col11[15];
   result_col11[17] <= result_col11[16];
   result_col11[18] <= result_col11[17];
   result_col11[19] <= result_col11[18];
   result_col11[20] <= result_col11[19];
   result_col11[21] <= result_col11[20];
   result_col11[22] <= result_col11[21];
   result_col11[23] <= result_col11[22];
   result_col11[24] <= result_col11[23];
   result_col11[25] <= result_col11[24];
   result_col11[26] <= result_col11[25];
   result_col11[27] <= result_col11[26];
   result_col11[28] <= result_col11[27];
   result_col11[29] <= result_col11[28];
   result_col11[30] <= result_col11[29];
   result_col11[31] <= result_col11[30];
   result_col11[32] <= result_col11[31];
   result_col11[33] <= result_col11[32];
   result_col11[34] <= result_col11[33];
   result_col11[35] <= result_col11[34];
   result_col11[36] <= result_col11[35];
   result_col11[37] <= result_col11[36];
   result_col11[38] <= result_col11[37];
   result_col11[39] <= result_col11[38];
   result_col11[40] <= result_col11[39];
   result_col11[41] <= result_col11[40];
   result_col11[42] <= result_col11[41];
   result_col11[43] <= result_col11[42];
   result_col11[44] <= result_col11[43];
   result_col11[45] <= result_col11[44];
   result_col11[46] <= result_col11[45];
   result_col11[47] <= result_col11[46];
   result_col11[48] <= result_col11[47];
   result_col11[49] <= result_col11[48];
   result_col11[50] <= result_col11[49];
   result_col11[51] <= result_col11[50];
   result_col11[52] <= result_col11[51];
   result_col11[53] <= result_col11[52];
   result_col11[54] <= result_col11[53];
   result_col11[55] <= result_col11[54];
   result_col11[56] <= result_col11[55];
   result_col11[57] <= result_col11[56];
   result_col11[58] <= result_col11[57];
   result_col11[59] <= result_col11[58];
   result_col11[60] <= result_col11[59];
   result_col11[61] <= result_col11[60];
   result_col11[62] <= result_col11[61];
   result_col11[63] <= result_col11[62];
   result_col11[64] <= result_col11[63];
   result_col11[65] <= result_col11[64];
   result_col11[66] <= result_col11[65];
   result_col11[67] <= result_col11[66];
   result_col11[68] <= result_col11[67];
   result_col11[69] <= result_col11[68];
   result_col11[70] <= result_col11[69];
   result_col11[71] <= result_col11[70];
   result_col11[72] <= result_col11[71];
   result_col11[73] <= result_col11[72];
   result_col11[74] <= result_col11[73];
   result_col11[75] <= result_col11[74];
   result_col11[76] <= result_col11[75];
   result_col11[77] <= result_col11[76];
   result_col11[78] <= result_col11[77];
   result_col11[79] <= result_col11[78];
   result_col11[80] <= result_col11[79];
   result_col11[81] <= result_col11[80];
   result_col11[82] <= result_col11[81];
   result_col11[83] <= result_col11[82];
   result_col11[84] <= result_col11[83];
   result_col11[85] <= result_col11[84];
   result_col11[86] <= result_col11[85];
   result_col11[87] <= result_col11[86];
   result_col11[88] <= result_col11[87];
   result_col11[89] <= result_col11[88];
   result_col11[90] <= result_col11[89];
   result_col11[91] <= result_col11[90];
   result_col11[92] <= result_col11[91];
   result_col11[93] <= result_col11[92];
   result_col11[94] <= result_col11[93];
   result_col11[95] <= result_col11[94];
   result_col11[96] <= result_col11[95];
   result_col11[97] <= result_col11[96];
   result_col11[98] <= result_col11[97];
   result_col11[99] <= result_col11[98];
   result_col11[100] <= result_col11[99];
   result_col11[101] <= result_col11[100];
   result_col11[102] <= result_col11[101];
   result_col11[103] <= result_col11[102];
   result_col11[104] <= result_col11[103];
   result_col11[105] <= result_col11[104];
   result_col11[106] <= result_col11[105];
   result_col11[107] <= result_col11[106];
   result_col11[108] <= result_col11[107];
   result_col11[109] <= result_col11[108];
   result_col11[110] <= result_col11[109];
   result_col11[111] <= result_col11[110];
   result_col11[112] <= result_col11[111];
   result_col11[113] <= result_col11[112];
   result_col11[114] <= result_col11[113];
   result_col11[115] <= result_col11[114];
   result_col11[116] <= result_col11[115];
   result_col11[117] <= result_col11[116];
   result_col11[118] <= result_col11[117];
   result_col11[119] <= result_col11[118];
   result_col11[120] <= result_col11[119];
   result_col11[121] <= result_col11[120];
   result_col11[122] <= result_col11[121];
   result_col11[123] <= result_col11[122];
   result_col11[124] <= result_col11[123];
   result_col11[125] <= result_col11[124];
   result_col11[126] <= result_col11[125];
   result_col11[127] <= result_col11[126];
   result_col11[128] <= result_col11[127];
   result_col11[129] <= result_col11[128];
   result_col11[130] <= result_col11[129];
   result_col11[131] <= result_col11[130];
   result_col11[132] <= result_col11[131];
   result_col11[133] <= result_col11[132];
   result_col11[134] <= result_col11[133];
   result_col11[135] <= result_col11[134];
   result_col11[136] <= result_col11[135];
   result_col11[137] <= result_col11[136];
   result_col11[138] <= result_col11[137];
   result_col11[139] <= result_col11[138];
   result_col11[140] <= result_col11[139];
   result_col11[141] <= result_col11[140];
   result_col11[142] <= result_col11[141];
   result_col11[143] <= result_col11[142];
   result_col11[144] <= result_col11[143];
   result_col11[145] <= result_col11[144];
   result_col11[146] <= result_col11[145];
   result_col11[147] <= result_col11[146];
   result_col11[148] <= result_col11[147];
   result_col11[149] <= result_col11[148];
   result_col11[150] <= result_col11[149];
   result_col11[151] <= result_col11[150];
   result_col11[152] <= result_col11[151];
   result_col11[153] <= result_col11[152];
   result_col11[154] <= result_col11[153];
   result_col11[155] <= result_col11[154];

   result_col12[1] <= data_out_4_12;
   result_col12[2] <= result_col12[1];
   result_col12[3] <= result_col12[2];
   result_col12[4] <= result_col12[3];
   result_col12[5] <= result_col12[4];
   result_col12[6] <= result_col12[5];
   result_col12[7] <= result_col12[6];
   result_col12[8] <= result_col12[7];
   result_col12[9] <= result_col12[8];
   result_col12[10] <= result_col12[9];
   result_col12[11] <= result_col12[10];
   result_col12[12] <= result_col12[11];
   result_col12[13] <= result_col12[12];
   result_col12[14] <= result_col12[13];
   result_col12[15] <= result_col12[14];
   result_col12[16] <= result_col12[15];
   result_col12[17] <= result_col12[16];
   result_col12[18] <= result_col12[17];
   result_col12[19] <= result_col12[18];
   result_col12[20] <= result_col12[19];
   result_col12[21] <= result_col12[20];
   result_col12[22] <= result_col12[21];
   result_col12[23] <= result_col12[22];
   result_col12[24] <= result_col12[23];
   result_col12[25] <= result_col12[24];
   result_col12[26] <= result_col12[25];
   result_col12[27] <= result_col12[26];
   result_col12[28] <= result_col12[27];
   result_col12[29] <= result_col12[28];
   result_col12[30] <= result_col12[29];
   result_col12[31] <= result_col12[30];
   result_col12[32] <= result_col12[31];
   result_col12[33] <= result_col12[32];
   result_col12[34] <= result_col12[33];
   result_col12[35] <= result_col12[34];
   result_col12[36] <= result_col12[35];
   result_col12[37] <= result_col12[36];
   result_col12[38] <= result_col12[37];
   result_col12[39] <= result_col12[38];
   result_col12[40] <= result_col12[39];
   result_col12[41] <= result_col12[40];
   result_col12[42] <= result_col12[41];
   result_col12[43] <= result_col12[42];
   result_col12[44] <= result_col12[43];
   result_col12[45] <= result_col12[44];
   result_col12[46] <= result_col12[45];
   result_col12[47] <= result_col12[46];
   result_col12[48] <= result_col12[47];
   result_col12[49] <= result_col12[48];
   result_col12[50] <= result_col12[49];
   result_col12[51] <= result_col12[50];
   result_col12[52] <= result_col12[51];
   result_col12[53] <= result_col12[52];
   result_col12[54] <= result_col12[53];
   result_col12[55] <= result_col12[54];
   result_col12[56] <= result_col12[55];
   result_col12[57] <= result_col12[56];
   result_col12[58] <= result_col12[57];
   result_col12[59] <= result_col12[58];
   result_col12[60] <= result_col12[59];
   result_col12[61] <= result_col12[60];
   result_col12[62] <= result_col12[61];
   result_col12[63] <= result_col12[62];
   result_col12[64] <= result_col12[63];
   result_col12[65] <= result_col12[64];
   result_col12[66] <= result_col12[65];
   result_col12[67] <= result_col12[66];
   result_col12[68] <= result_col12[67];
   result_col12[69] <= result_col12[68];
   result_col12[70] <= result_col12[69];
   result_col12[71] <= result_col12[70];
   result_col12[72] <= result_col12[71];
   result_col12[73] <= result_col12[72];
   result_col12[74] <= result_col12[73];
   result_col12[75] <= result_col12[74];
   result_col12[76] <= result_col12[75];
   result_col12[77] <= result_col12[76];
   result_col12[78] <= result_col12[77];
   result_col12[79] <= result_col12[78];
   result_col12[80] <= result_col12[79];
   result_col12[81] <= result_col12[80];
   result_col12[82] <= result_col12[81];
   result_col12[83] <= result_col12[82];
   result_col12[84] <= result_col12[83];
   result_col12[85] <= result_col12[84];
   result_col12[86] <= result_col12[85];
   result_col12[87] <= result_col12[86];
   result_col12[88] <= result_col12[87];
   result_col12[89] <= result_col12[88];
   result_col12[90] <= result_col12[89];
   result_col12[91] <= result_col12[90];
   result_col12[92] <= result_col12[91];
   result_col12[93] <= result_col12[92];
   result_col12[94] <= result_col12[93];
   result_col12[95] <= result_col12[94];
   result_col12[96] <= result_col12[95];
   result_col12[97] <= result_col12[96];
   result_col12[98] <= result_col12[97];
   result_col12[99] <= result_col12[98];
   result_col12[100] <= result_col12[99];
   result_col12[101] <= result_col12[100];
   result_col12[102] <= result_col12[101];
   result_col12[103] <= result_col12[102];
   result_col12[104] <= result_col12[103];
   result_col12[105] <= result_col12[104];
   result_col12[106] <= result_col12[105];
   result_col12[107] <= result_col12[106];
   result_col12[108] <= result_col12[107];
   result_col12[109] <= result_col12[108];
   result_col12[110] <= result_col12[109];
   result_col12[111] <= result_col12[110];
   result_col12[112] <= result_col12[111];
   result_col12[113] <= result_col12[112];
   result_col12[114] <= result_col12[113];
   result_col12[115] <= result_col12[114];
   result_col12[116] <= result_col12[115];
   result_col12[117] <= result_col12[116];
   result_col12[118] <= result_col12[117];
   result_col12[119] <= result_col12[118];
   result_col12[120] <= result_col12[119];
   result_col12[121] <= result_col12[120];
   result_col12[122] <= result_col12[121];
   result_col12[123] <= result_col12[122];
   result_col12[124] <= result_col12[123];
   result_col12[125] <= result_col12[124];
   result_col12[126] <= result_col12[125];
   result_col12[127] <= result_col12[126];
   result_col12[128] <= result_col12[127];
   result_col12[129] <= result_col12[128];
   result_col12[130] <= result_col12[129];
   result_col12[131] <= result_col12[130];
   result_col12[132] <= result_col12[131];
   result_col12[133] <= result_col12[132];
   result_col12[134] <= result_col12[133];
   result_col12[135] <= result_col12[134];
   result_col12[136] <= result_col12[135];
   result_col12[137] <= result_col12[136];
   result_col12[138] <= result_col12[137];
   result_col12[139] <= result_col12[138];
   result_col12[140] <= result_col12[139];
   result_col12[141] <= result_col12[140];
   result_col12[142] <= result_col12[141];
   result_col12[143] <= result_col12[142];
   result_col12[144] <= result_col12[143];
   result_col12[145] <= result_col12[144];
   result_col12[146] <= result_col12[145];
   result_col12[147] <= result_col12[146];
   result_col12[148] <= result_col12[147];
   result_col12[149] <= result_col12[148];
   result_col12[150] <= result_col12[149];
   result_col12[151] <= result_col12[150];
   result_col12[152] <= result_col12[151];
   result_col12[153] <= result_col12[152];
   result_col12[154] <= result_col12[153];

   result_col13[1] <= data_out_4_13;
   result_col13[2] <= result_col13[1];
   result_col13[3] <= result_col13[2];
   result_col13[4] <= result_col13[3];
   result_col13[5] <= result_col13[4];
   result_col13[6] <= result_col13[5];
   result_col13[7] <= result_col13[6];
   result_col13[8] <= result_col13[7];
   result_col13[9] <= result_col13[8];
   result_col13[10] <= result_col13[9];
   result_col13[11] <= result_col13[10];
   result_col13[12] <= result_col13[11];
   result_col13[13] <= result_col13[12];
   result_col13[14] <= result_col13[13];
   result_col13[15] <= result_col13[14];
   result_col13[16] <= result_col13[15];
   result_col13[17] <= result_col13[16];
   result_col13[18] <= result_col13[17];
   result_col13[19] <= result_col13[18];
   result_col13[20] <= result_col13[19];
   result_col13[21] <= result_col13[20];
   result_col13[22] <= result_col13[21];
   result_col13[23] <= result_col13[22];
   result_col13[24] <= result_col13[23];
   result_col13[25] <= result_col13[24];
   result_col13[26] <= result_col13[25];
   result_col13[27] <= result_col13[26];
   result_col13[28] <= result_col13[27];
   result_col13[29] <= result_col13[28];
   result_col13[30] <= result_col13[29];
   result_col13[31] <= result_col13[30];
   result_col13[32] <= result_col13[31];
   result_col13[33] <= result_col13[32];
   result_col13[34] <= result_col13[33];
   result_col13[35] <= result_col13[34];
   result_col13[36] <= result_col13[35];
   result_col13[37] <= result_col13[36];
   result_col13[38] <= result_col13[37];
   result_col13[39] <= result_col13[38];
   result_col13[40] <= result_col13[39];
   result_col13[41] <= result_col13[40];
   result_col13[42] <= result_col13[41];
   result_col13[43] <= result_col13[42];
   result_col13[44] <= result_col13[43];
   result_col13[45] <= result_col13[44];
   result_col13[46] <= result_col13[45];
   result_col13[47] <= result_col13[46];
   result_col13[48] <= result_col13[47];
   result_col13[49] <= result_col13[48];
   result_col13[50] <= result_col13[49];
   result_col13[51] <= result_col13[50];
   result_col13[52] <= result_col13[51];
   result_col13[53] <= result_col13[52];
   result_col13[54] <= result_col13[53];
   result_col13[55] <= result_col13[54];
   result_col13[56] <= result_col13[55];
   result_col13[57] <= result_col13[56];
   result_col13[58] <= result_col13[57];
   result_col13[59] <= result_col13[58];
   result_col13[60] <= result_col13[59];
   result_col13[61] <= result_col13[60];
   result_col13[62] <= result_col13[61];
   result_col13[63] <= result_col13[62];
   result_col13[64] <= result_col13[63];
   result_col13[65] <= result_col13[64];
   result_col13[66] <= result_col13[65];
   result_col13[67] <= result_col13[66];
   result_col13[68] <= result_col13[67];
   result_col13[69] <= result_col13[68];
   result_col13[70] <= result_col13[69];
   result_col13[71] <= result_col13[70];
   result_col13[72] <= result_col13[71];
   result_col13[73] <= result_col13[72];
   result_col13[74] <= result_col13[73];
   result_col13[75] <= result_col13[74];
   result_col13[76] <= result_col13[75];
   result_col13[77] <= result_col13[76];
   result_col13[78] <= result_col13[77];
   result_col13[79] <= result_col13[78];
   result_col13[80] <= result_col13[79];
   result_col13[81] <= result_col13[80];
   result_col13[82] <= result_col13[81];
   result_col13[83] <= result_col13[82];
   result_col13[84] <= result_col13[83];
   result_col13[85] <= result_col13[84];
   result_col13[86] <= result_col13[85];
   result_col13[87] <= result_col13[86];
   result_col13[88] <= result_col13[87];
   result_col13[89] <= result_col13[88];
   result_col13[90] <= result_col13[89];
   result_col13[91] <= result_col13[90];
   result_col13[92] <= result_col13[91];
   result_col13[93] <= result_col13[92];
   result_col13[94] <= result_col13[93];
   result_col13[95] <= result_col13[94];
   result_col13[96] <= result_col13[95];
   result_col13[97] <= result_col13[96];
   result_col13[98] <= result_col13[97];
   result_col13[99] <= result_col13[98];
   result_col13[100] <= result_col13[99];
   result_col13[101] <= result_col13[100];
   result_col13[102] <= result_col13[101];
   result_col13[103] <= result_col13[102];
   result_col13[104] <= result_col13[103];
   result_col13[105] <= result_col13[104];
   result_col13[106] <= result_col13[105];
   result_col13[107] <= result_col13[106];
   result_col13[108] <= result_col13[107];
   result_col13[109] <= result_col13[108];
   result_col13[110] <= result_col13[109];
   result_col13[111] <= result_col13[110];
   result_col13[112] <= result_col13[111];
   result_col13[113] <= result_col13[112];
   result_col13[114] <= result_col13[113];
   result_col13[115] <= result_col13[114];
   result_col13[116] <= result_col13[115];
   result_col13[117] <= result_col13[116];
   result_col13[118] <= result_col13[117];
   result_col13[119] <= result_col13[118];
   result_col13[120] <= result_col13[119];
   result_col13[121] <= result_col13[120];
   result_col13[122] <= result_col13[121];
   result_col13[123] <= result_col13[122];
   result_col13[124] <= result_col13[123];
   result_col13[125] <= result_col13[124];
   result_col13[126] <= result_col13[125];
   result_col13[127] <= result_col13[126];
   result_col13[128] <= result_col13[127];
   result_col13[129] <= result_col13[128];
   result_col13[130] <= result_col13[129];
   result_col13[131] <= result_col13[130];
   result_col13[132] <= result_col13[131];
   result_col13[133] <= result_col13[132];
   result_col13[134] <= result_col13[133];
   result_col13[135] <= result_col13[134];
   result_col13[136] <= result_col13[135];
   result_col13[137] <= result_col13[136];
   result_col13[138] <= result_col13[137];
   result_col13[139] <= result_col13[138];
   result_col13[140] <= result_col13[139];
   result_col13[141] <= result_col13[140];
   result_col13[142] <= result_col13[141];
   result_col13[143] <= result_col13[142];
   result_col13[144] <= result_col13[143];
   result_col13[145] <= result_col13[144];
   result_col13[146] <= result_col13[145];
   result_col13[147] <= result_col13[146];
   result_col13[148] <= result_col13[147];
   result_col13[149] <= result_col13[148];
   result_col13[150] <= result_col13[149];
   result_col13[151] <= result_col13[150];
   result_col13[152] <= result_col13[151];
   result_col13[153] <= result_col13[152];

   result_col14[1] <= data_out_4_14;
   result_col14[2] <= result_col14[1];
   result_col14[3] <= result_col14[2];
   result_col14[4] <= result_col14[3];
   result_col14[5] <= result_col14[4];
   result_col14[6] <= result_col14[5];
   result_col14[7] <= result_col14[6];
   result_col14[8] <= result_col14[7];
   result_col14[9] <= result_col14[8];
   result_col14[10] <= result_col14[9];
   result_col14[11] <= result_col14[10];
   result_col14[12] <= result_col14[11];
   result_col14[13] <= result_col14[12];
   result_col14[14] <= result_col14[13];
   result_col14[15] <= result_col14[14];
   result_col14[16] <= result_col14[15];
   result_col14[17] <= result_col14[16];
   result_col14[18] <= result_col14[17];
   result_col14[19] <= result_col14[18];
   result_col14[20] <= result_col14[19];
   result_col14[21] <= result_col14[20];
   result_col14[22] <= result_col14[21];
   result_col14[23] <= result_col14[22];
   result_col14[24] <= result_col14[23];
   result_col14[25] <= result_col14[24];
   result_col14[26] <= result_col14[25];
   result_col14[27] <= result_col14[26];
   result_col14[28] <= result_col14[27];
   result_col14[29] <= result_col14[28];
   result_col14[30] <= result_col14[29];
   result_col14[31] <= result_col14[30];
   result_col14[32] <= result_col14[31];
   result_col14[33] <= result_col14[32];
   result_col14[34] <= result_col14[33];
   result_col14[35] <= result_col14[34];
   result_col14[36] <= result_col14[35];
   result_col14[37] <= result_col14[36];
   result_col14[38] <= result_col14[37];
   result_col14[39] <= result_col14[38];
   result_col14[40] <= result_col14[39];
   result_col14[41] <= result_col14[40];
   result_col14[42] <= result_col14[41];
   result_col14[43] <= result_col14[42];
   result_col14[44] <= result_col14[43];
   result_col14[45] <= result_col14[44];
   result_col14[46] <= result_col14[45];
   result_col14[47] <= result_col14[46];
   result_col14[48] <= result_col14[47];
   result_col14[49] <= result_col14[48];
   result_col14[50] <= result_col14[49];
   result_col14[51] <= result_col14[50];
   result_col14[52] <= result_col14[51];
   result_col14[53] <= result_col14[52];
   result_col14[54] <= result_col14[53];
   result_col14[55] <= result_col14[54];
   result_col14[56] <= result_col14[55];
   result_col14[57] <= result_col14[56];
   result_col14[58] <= result_col14[57];
   result_col14[59] <= result_col14[58];
   result_col14[60] <= result_col14[59];
   result_col14[61] <= result_col14[60];
   result_col14[62] <= result_col14[61];
   result_col14[63] <= result_col14[62];
   result_col14[64] <= result_col14[63];
   result_col14[65] <= result_col14[64];
   result_col14[66] <= result_col14[65];
   result_col14[67] <= result_col14[66];
   result_col14[68] <= result_col14[67];
   result_col14[69] <= result_col14[68];
   result_col14[70] <= result_col14[69];
   result_col14[71] <= result_col14[70];
   result_col14[72] <= result_col14[71];
   result_col14[73] <= result_col14[72];
   result_col14[74] <= result_col14[73];
   result_col14[75] <= result_col14[74];
   result_col14[76] <= result_col14[75];
   result_col14[77] <= result_col14[76];
   result_col14[78] <= result_col14[77];
   result_col14[79] <= result_col14[78];
   result_col14[80] <= result_col14[79];
   result_col14[81] <= result_col14[80];
   result_col14[82] <= result_col14[81];
   result_col14[83] <= result_col14[82];
   result_col14[84] <= result_col14[83];
   result_col14[85] <= result_col14[84];
   result_col14[86] <= result_col14[85];
   result_col14[87] <= result_col14[86];
   result_col14[88] <= result_col14[87];
   result_col14[89] <= result_col14[88];
   result_col14[90] <= result_col14[89];
   result_col14[91] <= result_col14[90];
   result_col14[92] <= result_col14[91];
   result_col14[93] <= result_col14[92];
   result_col14[94] <= result_col14[93];
   result_col14[95] <= result_col14[94];
   result_col14[96] <= result_col14[95];
   result_col14[97] <= result_col14[96];
   result_col14[98] <= result_col14[97];
   result_col14[99] <= result_col14[98];
   result_col14[100] <= result_col14[99];
   result_col14[101] <= result_col14[100];
   result_col14[102] <= result_col14[101];
   result_col14[103] <= result_col14[102];
   result_col14[104] <= result_col14[103];
   result_col14[105] <= result_col14[104];
   result_col14[106] <= result_col14[105];
   result_col14[107] <= result_col14[106];
   result_col14[108] <= result_col14[107];
   result_col14[109] <= result_col14[108];
   result_col14[110] <= result_col14[109];
   result_col14[111] <= result_col14[110];
   result_col14[112] <= result_col14[111];
   result_col14[113] <= result_col14[112];
   result_col14[114] <= result_col14[113];
   result_col14[115] <= result_col14[114];
   result_col14[116] <= result_col14[115];
   result_col14[117] <= result_col14[116];
   result_col14[118] <= result_col14[117];
   result_col14[119] <= result_col14[118];
   result_col14[120] <= result_col14[119];
   result_col14[121] <= result_col14[120];
   result_col14[122] <= result_col14[121];
   result_col14[123] <= result_col14[122];
   result_col14[124] <= result_col14[123];
   result_col14[125] <= result_col14[124];
   result_col14[126] <= result_col14[125];
   result_col14[127] <= result_col14[126];
   result_col14[128] <= result_col14[127];
   result_col14[129] <= result_col14[128];
   result_col14[130] <= result_col14[129];
   result_col14[131] <= result_col14[130];
   result_col14[132] <= result_col14[131];
   result_col14[133] <= result_col14[132];
   result_col14[134] <= result_col14[133];
   result_col14[135] <= result_col14[134];
   result_col14[136] <= result_col14[135];
   result_col14[137] <= result_col14[136];
   result_col14[138] <= result_col14[137];
   result_col14[139] <= result_col14[138];
   result_col14[140] <= result_col14[139];
   result_col14[141] <= result_col14[140];
   result_col14[142] <= result_col14[141];
   result_col14[143] <= result_col14[142];
   result_col14[144] <= result_col14[143];
   result_col14[145] <= result_col14[144];
   result_col14[146] <= result_col14[145];
   result_col14[147] <= result_col14[146];
   result_col14[148] <= result_col14[147];
   result_col14[149] <= result_col14[148];
   result_col14[150] <= result_col14[149];
   result_col14[151] <= result_col14[150];
   result_col14[152] <= result_col14[151];

   result_col15[1] <= data_out_4_15;
   result_col15[2] <= result_col15[1];
   result_col15[3] <= result_col15[2];
   result_col15[4] <= result_col15[3];
   result_col15[5] <= result_col15[4];
   result_col15[6] <= result_col15[5];
   result_col15[7] <= result_col15[6];
   result_col15[8] <= result_col15[7];
   result_col15[9] <= result_col15[8];
   result_col15[10] <= result_col15[9];
   result_col15[11] <= result_col15[10];
   result_col15[12] <= result_col15[11];
   result_col15[13] <= result_col15[12];
   result_col15[14] <= result_col15[13];
   result_col15[15] <= result_col15[14];
   result_col15[16] <= result_col15[15];
   result_col15[17] <= result_col15[16];
   result_col15[18] <= result_col15[17];
   result_col15[19] <= result_col15[18];
   result_col15[20] <= result_col15[19];
   result_col15[21] <= result_col15[20];
   result_col15[22] <= result_col15[21];
   result_col15[23] <= result_col15[22];
   result_col15[24] <= result_col15[23];
   result_col15[25] <= result_col15[24];
   result_col15[26] <= result_col15[25];
   result_col15[27] <= result_col15[26];
   result_col15[28] <= result_col15[27];
   result_col15[29] <= result_col15[28];
   result_col15[30] <= result_col15[29];
   result_col15[31] <= result_col15[30];
   result_col15[32] <= result_col15[31];
   result_col15[33] <= result_col15[32];
   result_col15[34] <= result_col15[33];
   result_col15[35] <= result_col15[34];
   result_col15[36] <= result_col15[35];
   result_col15[37] <= result_col15[36];
   result_col15[38] <= result_col15[37];
   result_col15[39] <= result_col15[38];
   result_col15[40] <= result_col15[39];
   result_col15[41] <= result_col15[40];
   result_col15[42] <= result_col15[41];
   result_col15[43] <= result_col15[42];
   result_col15[44] <= result_col15[43];
   result_col15[45] <= result_col15[44];
   result_col15[46] <= result_col15[45];
   result_col15[47] <= result_col15[46];
   result_col15[48] <= result_col15[47];
   result_col15[49] <= result_col15[48];
   result_col15[50] <= result_col15[49];
   result_col15[51] <= result_col15[50];
   result_col15[52] <= result_col15[51];
   result_col15[53] <= result_col15[52];
   result_col15[54] <= result_col15[53];
   result_col15[55] <= result_col15[54];
   result_col15[56] <= result_col15[55];
   result_col15[57] <= result_col15[56];
   result_col15[58] <= result_col15[57];
   result_col15[59] <= result_col15[58];
   result_col15[60] <= result_col15[59];
   result_col15[61] <= result_col15[60];
   result_col15[62] <= result_col15[61];
   result_col15[63] <= result_col15[62];
   result_col15[64] <= result_col15[63];
   result_col15[65] <= result_col15[64];
   result_col15[66] <= result_col15[65];
   result_col15[67] <= result_col15[66];
   result_col15[68] <= result_col15[67];
   result_col15[69] <= result_col15[68];
   result_col15[70] <= result_col15[69];
   result_col15[71] <= result_col15[70];
   result_col15[72] <= result_col15[71];
   result_col15[73] <= result_col15[72];
   result_col15[74] <= result_col15[73];
   result_col15[75] <= result_col15[74];
   result_col15[76] <= result_col15[75];
   result_col15[77] <= result_col15[76];
   result_col15[78] <= result_col15[77];
   result_col15[79] <= result_col15[78];
   result_col15[80] <= result_col15[79];
   result_col15[81] <= result_col15[80];
   result_col15[82] <= result_col15[81];
   result_col15[83] <= result_col15[82];
   result_col15[84] <= result_col15[83];
   result_col15[85] <= result_col15[84];
   result_col15[86] <= result_col15[85];
   result_col15[87] <= result_col15[86];
   result_col15[88] <= result_col15[87];
   result_col15[89] <= result_col15[88];
   result_col15[90] <= result_col15[89];
   result_col15[91] <= result_col15[90];
   result_col15[92] <= result_col15[91];
   result_col15[93] <= result_col15[92];
   result_col15[94] <= result_col15[93];
   result_col15[95] <= result_col15[94];
   result_col15[96] <= result_col15[95];
   result_col15[97] <= result_col15[96];
   result_col15[98] <= result_col15[97];
   result_col15[99] <= result_col15[98];
   result_col15[100] <= result_col15[99];
   result_col15[101] <= result_col15[100];
   result_col15[102] <= result_col15[101];
   result_col15[103] <= result_col15[102];
   result_col15[104] <= result_col15[103];
   result_col15[105] <= result_col15[104];
   result_col15[106] <= result_col15[105];
   result_col15[107] <= result_col15[106];
   result_col15[108] <= result_col15[107];
   result_col15[109] <= result_col15[108];
   result_col15[110] <= result_col15[109];
   result_col15[111] <= result_col15[110];
   result_col15[112] <= result_col15[111];
   result_col15[113] <= result_col15[112];
   result_col15[114] <= result_col15[113];
   result_col15[115] <= result_col15[114];
   result_col15[116] <= result_col15[115];
   result_col15[117] <= result_col15[116];
   result_col15[118] <= result_col15[117];
   result_col15[119] <= result_col15[118];
   result_col15[120] <= result_col15[119];
   result_col15[121] <= result_col15[120];
   result_col15[122] <= result_col15[121];
   result_col15[123] <= result_col15[122];
   result_col15[124] <= result_col15[123];
   result_col15[125] <= result_col15[124];
   result_col15[126] <= result_col15[125];
   result_col15[127] <= result_col15[126];
   result_col15[128] <= result_col15[127];
   result_col15[129] <= result_col15[128];
   result_col15[130] <= result_col15[129];
   result_col15[131] <= result_col15[130];
   result_col15[132] <= result_col15[131];
   result_col15[133] <= result_col15[132];
   result_col15[134] <= result_col15[133];
   result_col15[135] <= result_col15[134];
   result_col15[136] <= result_col15[135];
   result_col15[137] <= result_col15[136];
   result_col15[138] <= result_col15[137];
   result_col15[139] <= result_col15[138];
   result_col15[140] <= result_col15[139];
   result_col15[141] <= result_col15[140];
   result_col15[142] <= result_col15[141];
   result_col15[143] <= result_col15[142];
   result_col15[144] <= result_col15[143];
   result_col15[145] <= result_col15[144];
   result_col15[146] <= result_col15[145];
   result_col15[147] <= result_col15[146];
   result_col15[148] <= result_col15[147];
   result_col15[149] <= result_col15[148];
   result_col15[150] <= result_col15[149];
   result_col15[151] <= result_col15[150];

   result_col16[1] <= data_out_4_16;
   result_col16[2] <= result_col16[1];
   result_col16[3] <= result_col16[2];
   result_col16[4] <= result_col16[3];
   result_col16[5] <= result_col16[4];
   result_col16[6] <= result_col16[5];
   result_col16[7] <= result_col16[6];
   result_col16[8] <= result_col16[7];
   result_col16[9] <= result_col16[8];
   result_col16[10] <= result_col16[9];
   result_col16[11] <= result_col16[10];
   result_col16[12] <= result_col16[11];
   result_col16[13] <= result_col16[12];
   result_col16[14] <= result_col16[13];
   result_col16[15] <= result_col16[14];
   result_col16[16] <= result_col16[15];
   result_col16[17] <= result_col16[16];
   result_col16[18] <= result_col16[17];
   result_col16[19] <= result_col16[18];
   result_col16[20] <= result_col16[19];
   result_col16[21] <= result_col16[20];
   result_col16[22] <= result_col16[21];
   result_col16[23] <= result_col16[22];
   result_col16[24] <= result_col16[23];
   result_col16[25] <= result_col16[24];
   result_col16[26] <= result_col16[25];
   result_col16[27] <= result_col16[26];
   result_col16[28] <= result_col16[27];
   result_col16[29] <= result_col16[28];
   result_col16[30] <= result_col16[29];
   result_col16[31] <= result_col16[30];
   result_col16[32] <= result_col16[31];
   result_col16[33] <= result_col16[32];
   result_col16[34] <= result_col16[33];
   result_col16[35] <= result_col16[34];
   result_col16[36] <= result_col16[35];
   result_col16[37] <= result_col16[36];
   result_col16[38] <= result_col16[37];
   result_col16[39] <= result_col16[38];
   result_col16[40] <= result_col16[39];
   result_col16[41] <= result_col16[40];
   result_col16[42] <= result_col16[41];
   result_col16[43] <= result_col16[42];
   result_col16[44] <= result_col16[43];
   result_col16[45] <= result_col16[44];
   result_col16[46] <= result_col16[45];
   result_col16[47] <= result_col16[46];
   result_col16[48] <= result_col16[47];
   result_col16[49] <= result_col16[48];
   result_col16[50] <= result_col16[49];
   result_col16[51] <= result_col16[50];
   result_col16[52] <= result_col16[51];
   result_col16[53] <= result_col16[52];
   result_col16[54] <= result_col16[53];
   result_col16[55] <= result_col16[54];
   result_col16[56] <= result_col16[55];
   result_col16[57] <= result_col16[56];
   result_col16[58] <= result_col16[57];
   result_col16[59] <= result_col16[58];
   result_col16[60] <= result_col16[59];
   result_col16[61] <= result_col16[60];
   result_col16[62] <= result_col16[61];
   result_col16[63] <= result_col16[62];
   result_col16[64] <= result_col16[63];
   result_col16[65] <= result_col16[64];
   result_col16[66] <= result_col16[65];
   result_col16[67] <= result_col16[66];
   result_col16[68] <= result_col16[67];
   result_col16[69] <= result_col16[68];
   result_col16[70] <= result_col16[69];
   result_col16[71] <= result_col16[70];
   result_col16[72] <= result_col16[71];
   result_col16[73] <= result_col16[72];
   result_col16[74] <= result_col16[73];
   result_col16[75] <= result_col16[74];
   result_col16[76] <= result_col16[75];
   result_col16[77] <= result_col16[76];
   result_col16[78] <= result_col16[77];
   result_col16[79] <= result_col16[78];
   result_col16[80] <= result_col16[79];
   result_col16[81] <= result_col16[80];
   result_col16[82] <= result_col16[81];
   result_col16[83] <= result_col16[82];
   result_col16[84] <= result_col16[83];
   result_col16[85] <= result_col16[84];
   result_col16[86] <= result_col16[85];
   result_col16[87] <= result_col16[86];
   result_col16[88] <= result_col16[87];
   result_col16[89] <= result_col16[88];
   result_col16[90] <= result_col16[89];
   result_col16[91] <= result_col16[90];
   result_col16[92] <= result_col16[91];
   result_col16[93] <= result_col16[92];
   result_col16[94] <= result_col16[93];
   result_col16[95] <= result_col16[94];
   result_col16[96] <= result_col16[95];
   result_col16[97] <= result_col16[96];
   result_col16[98] <= result_col16[97];
   result_col16[99] <= result_col16[98];
   result_col16[100] <= result_col16[99];
   result_col16[101] <= result_col16[100];
   result_col16[102] <= result_col16[101];
   result_col16[103] <= result_col16[102];
   result_col16[104] <= result_col16[103];
   result_col16[105] <= result_col16[104];
   result_col16[106] <= result_col16[105];
   result_col16[107] <= result_col16[106];
   result_col16[108] <= result_col16[107];
   result_col16[109] <= result_col16[108];
   result_col16[110] <= result_col16[109];
   result_col16[111] <= result_col16[110];
   result_col16[112] <= result_col16[111];
   result_col16[113] <= result_col16[112];
   result_col16[114] <= result_col16[113];
   result_col16[115] <= result_col16[114];
   result_col16[116] <= result_col16[115];
   result_col16[117] <= result_col16[116];
   result_col16[118] <= result_col16[117];
   result_col16[119] <= result_col16[118];
   result_col16[120] <= result_col16[119];
   result_col16[121] <= result_col16[120];
   result_col16[122] <= result_col16[121];
   result_col16[123] <= result_col16[122];
   result_col16[124] <= result_col16[123];
   result_col16[125] <= result_col16[124];
   result_col16[126] <= result_col16[125];
   result_col16[127] <= result_col16[126];
   result_col16[128] <= result_col16[127];
   result_col16[129] <= result_col16[128];
   result_col16[130] <= result_col16[129];
   result_col16[131] <= result_col16[130];
   result_col16[132] <= result_col16[131];
   result_col16[133] <= result_col16[132];
   result_col16[134] <= result_col16[133];
   result_col16[135] <= result_col16[134];
   result_col16[136] <= result_col16[135];
   result_col16[137] <= result_col16[136];
   result_col16[138] <= result_col16[137];
   result_col16[139] <= result_col16[138];
   result_col16[140] <= result_col16[139];
   result_col16[141] <= result_col16[140];
   result_col16[142] <= result_col16[141];
   result_col16[143] <= result_col16[142];
   result_col16[144] <= result_col16[143];
   result_col16[145] <= result_col16[144];
   result_col16[146] <= result_col16[145];
   result_col16[147] <= result_col16[146];
   result_col16[148] <= result_col16[147];
   result_col16[149] <= result_col16[148];
   result_col16[150] <= result_col16[149];

   result_col17[1] <= data_out_4_17;
   result_col17[2] <= result_col17[1];
   result_col17[3] <= result_col17[2];
   result_col17[4] <= result_col17[3];
   result_col17[5] <= result_col17[4];
   result_col17[6] <= result_col17[5];
   result_col17[7] <= result_col17[6];
   result_col17[8] <= result_col17[7];
   result_col17[9] <= result_col17[8];
   result_col17[10] <= result_col17[9];
   result_col17[11] <= result_col17[10];
   result_col17[12] <= result_col17[11];
   result_col17[13] <= result_col17[12];
   result_col17[14] <= result_col17[13];
   result_col17[15] <= result_col17[14];
   result_col17[16] <= result_col17[15];
   result_col17[17] <= result_col17[16];
   result_col17[18] <= result_col17[17];
   result_col17[19] <= result_col17[18];
   result_col17[20] <= result_col17[19];
   result_col17[21] <= result_col17[20];
   result_col17[22] <= result_col17[21];
   result_col17[23] <= result_col17[22];
   result_col17[24] <= result_col17[23];
   result_col17[25] <= result_col17[24];
   result_col17[26] <= result_col17[25];
   result_col17[27] <= result_col17[26];
   result_col17[28] <= result_col17[27];
   result_col17[29] <= result_col17[28];
   result_col17[30] <= result_col17[29];
   result_col17[31] <= result_col17[30];
   result_col17[32] <= result_col17[31];
   result_col17[33] <= result_col17[32];
   result_col17[34] <= result_col17[33];
   result_col17[35] <= result_col17[34];
   result_col17[36] <= result_col17[35];
   result_col17[37] <= result_col17[36];
   result_col17[38] <= result_col17[37];
   result_col17[39] <= result_col17[38];
   result_col17[40] <= result_col17[39];
   result_col17[41] <= result_col17[40];
   result_col17[42] <= result_col17[41];
   result_col17[43] <= result_col17[42];
   result_col17[44] <= result_col17[43];
   result_col17[45] <= result_col17[44];
   result_col17[46] <= result_col17[45];
   result_col17[47] <= result_col17[46];
   result_col17[48] <= result_col17[47];
   result_col17[49] <= result_col17[48];
   result_col17[50] <= result_col17[49];
   result_col17[51] <= result_col17[50];
   result_col17[52] <= result_col17[51];
   result_col17[53] <= result_col17[52];
   result_col17[54] <= result_col17[53];
   result_col17[55] <= result_col17[54];
   result_col17[56] <= result_col17[55];
   result_col17[57] <= result_col17[56];
   result_col17[58] <= result_col17[57];
   result_col17[59] <= result_col17[58];
   result_col17[60] <= result_col17[59];
   result_col17[61] <= result_col17[60];
   result_col17[62] <= result_col17[61];
   result_col17[63] <= result_col17[62];
   result_col17[64] <= result_col17[63];
   result_col17[65] <= result_col17[64];
   result_col17[66] <= result_col17[65];
   result_col17[67] <= result_col17[66];
   result_col17[68] <= result_col17[67];
   result_col17[69] <= result_col17[68];
   result_col17[70] <= result_col17[69];
   result_col17[71] <= result_col17[70];
   result_col17[72] <= result_col17[71];
   result_col17[73] <= result_col17[72];
   result_col17[74] <= result_col17[73];
   result_col17[75] <= result_col17[74];
   result_col17[76] <= result_col17[75];
   result_col17[77] <= result_col17[76];
   result_col17[78] <= result_col17[77];
   result_col17[79] <= result_col17[78];
   result_col17[80] <= result_col17[79];
   result_col17[81] <= result_col17[80];
   result_col17[82] <= result_col17[81];
   result_col17[83] <= result_col17[82];
   result_col17[84] <= result_col17[83];
   result_col17[85] <= result_col17[84];
   result_col17[86] <= result_col17[85];
   result_col17[87] <= result_col17[86];
   result_col17[88] <= result_col17[87];
   result_col17[89] <= result_col17[88];
   result_col17[90] <= result_col17[89];
   result_col17[91] <= result_col17[90];
   result_col17[92] <= result_col17[91];
   result_col17[93] <= result_col17[92];
   result_col17[94] <= result_col17[93];
   result_col17[95] <= result_col17[94];
   result_col17[96] <= result_col17[95];
   result_col17[97] <= result_col17[96];
   result_col17[98] <= result_col17[97];
   result_col17[99] <= result_col17[98];
   result_col17[100] <= result_col17[99];
   result_col17[101] <= result_col17[100];
   result_col17[102] <= result_col17[101];
   result_col17[103] <= result_col17[102];
   result_col17[104] <= result_col17[103];
   result_col17[105] <= result_col17[104];
   result_col17[106] <= result_col17[105];
   result_col17[107] <= result_col17[106];
   result_col17[108] <= result_col17[107];
   result_col17[109] <= result_col17[108];
   result_col17[110] <= result_col17[109];
   result_col17[111] <= result_col17[110];
   result_col17[112] <= result_col17[111];
   result_col17[113] <= result_col17[112];
   result_col17[114] <= result_col17[113];
   result_col17[115] <= result_col17[114];
   result_col17[116] <= result_col17[115];
   result_col17[117] <= result_col17[116];
   result_col17[118] <= result_col17[117];
   result_col17[119] <= result_col17[118];
   result_col17[120] <= result_col17[119];
   result_col17[121] <= result_col17[120];
   result_col17[122] <= result_col17[121];
   result_col17[123] <= result_col17[122];
   result_col17[124] <= result_col17[123];
   result_col17[125] <= result_col17[124];
   result_col17[126] <= result_col17[125];
   result_col17[127] <= result_col17[126];
   result_col17[128] <= result_col17[127];
   result_col17[129] <= result_col17[128];
   result_col17[130] <= result_col17[129];
   result_col17[131] <= result_col17[130];
   result_col17[132] <= result_col17[131];
   result_col17[133] <= result_col17[132];
   result_col17[134] <= result_col17[133];
   result_col17[135] <= result_col17[134];
   result_col17[136] <= result_col17[135];
   result_col17[137] <= result_col17[136];
   result_col17[138] <= result_col17[137];
   result_col17[139] <= result_col17[138];
   result_col17[140] <= result_col17[139];
   result_col17[141] <= result_col17[140];
   result_col17[142] <= result_col17[141];
   result_col17[143] <= result_col17[142];
   result_col17[144] <= result_col17[143];
   result_col17[145] <= result_col17[144];
   result_col17[146] <= result_col17[145];
   result_col17[147] <= result_col17[146];
   result_col17[148] <= result_col17[147];
   result_col17[149] <= result_col17[148];

   result_col18[1] <= data_out_4_18;
   result_col18[2] <= result_col18[1];
   result_col18[3] <= result_col18[2];
   result_col18[4] <= result_col18[3];
   result_col18[5] <= result_col18[4];
   result_col18[6] <= result_col18[5];
   result_col18[7] <= result_col18[6];
   result_col18[8] <= result_col18[7];
   result_col18[9] <= result_col18[8];
   result_col18[10] <= result_col18[9];
   result_col18[11] <= result_col18[10];
   result_col18[12] <= result_col18[11];
   result_col18[13] <= result_col18[12];
   result_col18[14] <= result_col18[13];
   result_col18[15] <= result_col18[14];
   result_col18[16] <= result_col18[15];
   result_col18[17] <= result_col18[16];
   result_col18[18] <= result_col18[17];
   result_col18[19] <= result_col18[18];
   result_col18[20] <= result_col18[19];
   result_col18[21] <= result_col18[20];
   result_col18[22] <= result_col18[21];
   result_col18[23] <= result_col18[22];
   result_col18[24] <= result_col18[23];
   result_col18[25] <= result_col18[24];
   result_col18[26] <= result_col18[25];
   result_col18[27] <= result_col18[26];
   result_col18[28] <= result_col18[27];
   result_col18[29] <= result_col18[28];
   result_col18[30] <= result_col18[29];
   result_col18[31] <= result_col18[30];
   result_col18[32] <= result_col18[31];
   result_col18[33] <= result_col18[32];
   result_col18[34] <= result_col18[33];
   result_col18[35] <= result_col18[34];
   result_col18[36] <= result_col18[35];
   result_col18[37] <= result_col18[36];
   result_col18[38] <= result_col18[37];
   result_col18[39] <= result_col18[38];
   result_col18[40] <= result_col18[39];
   result_col18[41] <= result_col18[40];
   result_col18[42] <= result_col18[41];
   result_col18[43] <= result_col18[42];
   result_col18[44] <= result_col18[43];
   result_col18[45] <= result_col18[44];
   result_col18[46] <= result_col18[45];
   result_col18[47] <= result_col18[46];
   result_col18[48] <= result_col18[47];
   result_col18[49] <= result_col18[48];
   result_col18[50] <= result_col18[49];
   result_col18[51] <= result_col18[50];
   result_col18[52] <= result_col18[51];
   result_col18[53] <= result_col18[52];
   result_col18[54] <= result_col18[53];
   result_col18[55] <= result_col18[54];
   result_col18[56] <= result_col18[55];
   result_col18[57] <= result_col18[56];
   result_col18[58] <= result_col18[57];
   result_col18[59] <= result_col18[58];
   result_col18[60] <= result_col18[59];
   result_col18[61] <= result_col18[60];
   result_col18[62] <= result_col18[61];
   result_col18[63] <= result_col18[62];
   result_col18[64] <= result_col18[63];
   result_col18[65] <= result_col18[64];
   result_col18[66] <= result_col18[65];
   result_col18[67] <= result_col18[66];
   result_col18[68] <= result_col18[67];
   result_col18[69] <= result_col18[68];
   result_col18[70] <= result_col18[69];
   result_col18[71] <= result_col18[70];
   result_col18[72] <= result_col18[71];
   result_col18[73] <= result_col18[72];
   result_col18[74] <= result_col18[73];
   result_col18[75] <= result_col18[74];
   result_col18[76] <= result_col18[75];
   result_col18[77] <= result_col18[76];
   result_col18[78] <= result_col18[77];
   result_col18[79] <= result_col18[78];
   result_col18[80] <= result_col18[79];
   result_col18[81] <= result_col18[80];
   result_col18[82] <= result_col18[81];
   result_col18[83] <= result_col18[82];
   result_col18[84] <= result_col18[83];
   result_col18[85] <= result_col18[84];
   result_col18[86] <= result_col18[85];
   result_col18[87] <= result_col18[86];
   result_col18[88] <= result_col18[87];
   result_col18[89] <= result_col18[88];
   result_col18[90] <= result_col18[89];
   result_col18[91] <= result_col18[90];
   result_col18[92] <= result_col18[91];
   result_col18[93] <= result_col18[92];
   result_col18[94] <= result_col18[93];
   result_col18[95] <= result_col18[94];
   result_col18[96] <= result_col18[95];
   result_col18[97] <= result_col18[96];
   result_col18[98] <= result_col18[97];
   result_col18[99] <= result_col18[98];
   result_col18[100] <= result_col18[99];
   result_col18[101] <= result_col18[100];
   result_col18[102] <= result_col18[101];
   result_col18[103] <= result_col18[102];
   result_col18[104] <= result_col18[103];
   result_col18[105] <= result_col18[104];
   result_col18[106] <= result_col18[105];
   result_col18[107] <= result_col18[106];
   result_col18[108] <= result_col18[107];
   result_col18[109] <= result_col18[108];
   result_col18[110] <= result_col18[109];
   result_col18[111] <= result_col18[110];
   result_col18[112] <= result_col18[111];
   result_col18[113] <= result_col18[112];
   result_col18[114] <= result_col18[113];
   result_col18[115] <= result_col18[114];
   result_col18[116] <= result_col18[115];
   result_col18[117] <= result_col18[116];
   result_col18[118] <= result_col18[117];
   result_col18[119] <= result_col18[118];
   result_col18[120] <= result_col18[119];
   result_col18[121] <= result_col18[120];
   result_col18[122] <= result_col18[121];
   result_col18[123] <= result_col18[122];
   result_col18[124] <= result_col18[123];
   result_col18[125] <= result_col18[124];
   result_col18[126] <= result_col18[125];
   result_col18[127] <= result_col18[126];
   result_col18[128] <= result_col18[127];
   result_col18[129] <= result_col18[128];
   result_col18[130] <= result_col18[129];
   result_col18[131] <= result_col18[130];
   result_col18[132] <= result_col18[131];
   result_col18[133] <= result_col18[132];
   result_col18[134] <= result_col18[133];
   result_col18[135] <= result_col18[134];
   result_col18[136] <= result_col18[135];
   result_col18[137] <= result_col18[136];
   result_col18[138] <= result_col18[137];
   result_col18[139] <= result_col18[138];
   result_col18[140] <= result_col18[139];
   result_col18[141] <= result_col18[140];
   result_col18[142] <= result_col18[141];
   result_col18[143] <= result_col18[142];
   result_col18[144] <= result_col18[143];
   result_col18[145] <= result_col18[144];
   result_col18[146] <= result_col18[145];
   result_col18[147] <= result_col18[146];
   result_col18[148] <= result_col18[147];

   result_col19[1] <= data_out_4_19;
   result_col19[2] <= result_col19[1];
   result_col19[3] <= result_col19[2];
   result_col19[4] <= result_col19[3];
   result_col19[5] <= result_col19[4];
   result_col19[6] <= result_col19[5];
   result_col19[7] <= result_col19[6];
   result_col19[8] <= result_col19[7];
   result_col19[9] <= result_col19[8];
   result_col19[10] <= result_col19[9];
   result_col19[11] <= result_col19[10];
   result_col19[12] <= result_col19[11];
   result_col19[13] <= result_col19[12];
   result_col19[14] <= result_col19[13];
   result_col19[15] <= result_col19[14];
   result_col19[16] <= result_col19[15];
   result_col19[17] <= result_col19[16];
   result_col19[18] <= result_col19[17];
   result_col19[19] <= result_col19[18];
   result_col19[20] <= result_col19[19];
   result_col19[21] <= result_col19[20];
   result_col19[22] <= result_col19[21];
   result_col19[23] <= result_col19[22];
   result_col19[24] <= result_col19[23];
   result_col19[25] <= result_col19[24];
   result_col19[26] <= result_col19[25];
   result_col19[27] <= result_col19[26];
   result_col19[28] <= result_col19[27];
   result_col19[29] <= result_col19[28];
   result_col19[30] <= result_col19[29];
   result_col19[31] <= result_col19[30];
   result_col19[32] <= result_col19[31];
   result_col19[33] <= result_col19[32];
   result_col19[34] <= result_col19[33];
   result_col19[35] <= result_col19[34];
   result_col19[36] <= result_col19[35];
   result_col19[37] <= result_col19[36];
   result_col19[38] <= result_col19[37];
   result_col19[39] <= result_col19[38];
   result_col19[40] <= result_col19[39];
   result_col19[41] <= result_col19[40];
   result_col19[42] <= result_col19[41];
   result_col19[43] <= result_col19[42];
   result_col19[44] <= result_col19[43];
   result_col19[45] <= result_col19[44];
   result_col19[46] <= result_col19[45];
   result_col19[47] <= result_col19[46];
   result_col19[48] <= result_col19[47];
   result_col19[49] <= result_col19[48];
   result_col19[50] <= result_col19[49];
   result_col19[51] <= result_col19[50];
   result_col19[52] <= result_col19[51];
   result_col19[53] <= result_col19[52];
   result_col19[54] <= result_col19[53];
   result_col19[55] <= result_col19[54];
   result_col19[56] <= result_col19[55];
   result_col19[57] <= result_col19[56];
   result_col19[58] <= result_col19[57];
   result_col19[59] <= result_col19[58];
   result_col19[60] <= result_col19[59];
   result_col19[61] <= result_col19[60];
   result_col19[62] <= result_col19[61];
   result_col19[63] <= result_col19[62];
   result_col19[64] <= result_col19[63];
   result_col19[65] <= result_col19[64];
   result_col19[66] <= result_col19[65];
   result_col19[67] <= result_col19[66];
   result_col19[68] <= result_col19[67];
   result_col19[69] <= result_col19[68];
   result_col19[70] <= result_col19[69];
   result_col19[71] <= result_col19[70];
   result_col19[72] <= result_col19[71];
   result_col19[73] <= result_col19[72];
   result_col19[74] <= result_col19[73];
   result_col19[75] <= result_col19[74];
   result_col19[76] <= result_col19[75];
   result_col19[77] <= result_col19[76];
   result_col19[78] <= result_col19[77];
   result_col19[79] <= result_col19[78];
   result_col19[80] <= result_col19[79];
   result_col19[81] <= result_col19[80];
   result_col19[82] <= result_col19[81];
   result_col19[83] <= result_col19[82];
   result_col19[84] <= result_col19[83];
   result_col19[85] <= result_col19[84];
   result_col19[86] <= result_col19[85];
   result_col19[87] <= result_col19[86];
   result_col19[88] <= result_col19[87];
   result_col19[89] <= result_col19[88];
   result_col19[90] <= result_col19[89];
   result_col19[91] <= result_col19[90];
   result_col19[92] <= result_col19[91];
   result_col19[93] <= result_col19[92];
   result_col19[94] <= result_col19[93];
   result_col19[95] <= result_col19[94];
   result_col19[96] <= result_col19[95];
   result_col19[97] <= result_col19[96];
   result_col19[98] <= result_col19[97];
   result_col19[99] <= result_col19[98];
   result_col19[100] <= result_col19[99];
   result_col19[101] <= result_col19[100];
   result_col19[102] <= result_col19[101];
   result_col19[103] <= result_col19[102];
   result_col19[104] <= result_col19[103];
   result_col19[105] <= result_col19[104];
   result_col19[106] <= result_col19[105];
   result_col19[107] <= result_col19[106];
   result_col19[108] <= result_col19[107];
   result_col19[109] <= result_col19[108];
   result_col19[110] <= result_col19[109];
   result_col19[111] <= result_col19[110];
   result_col19[112] <= result_col19[111];
   result_col19[113] <= result_col19[112];
   result_col19[114] <= result_col19[113];
   result_col19[115] <= result_col19[114];
   result_col19[116] <= result_col19[115];
   result_col19[117] <= result_col19[116];
   result_col19[118] <= result_col19[117];
   result_col19[119] <= result_col19[118];
   result_col19[120] <= result_col19[119];
   result_col19[121] <= result_col19[120];
   result_col19[122] <= result_col19[121];
   result_col19[123] <= result_col19[122];
   result_col19[124] <= result_col19[123];
   result_col19[125] <= result_col19[124];
   result_col19[126] <= result_col19[125];
   result_col19[127] <= result_col19[126];
   result_col19[128] <= result_col19[127];
   result_col19[129] <= result_col19[128];
   result_col19[130] <= result_col19[129];
   result_col19[131] <= result_col19[130];
   result_col19[132] <= result_col19[131];
   result_col19[133] <= result_col19[132];
   result_col19[134] <= result_col19[133];
   result_col19[135] <= result_col19[134];
   result_col19[136] <= result_col19[135];
   result_col19[137] <= result_col19[136];
   result_col19[138] <= result_col19[137];
   result_col19[139] <= result_col19[138];
   result_col19[140] <= result_col19[139];
   result_col19[141] <= result_col19[140];
   result_col19[142] <= result_col19[141];
   result_col19[143] <= result_col19[142];
   result_col19[144] <= result_col19[143];
   result_col19[145] <= result_col19[144];
   result_col19[146] <= result_col19[145];
   result_col19[147] <= result_col19[146];

   result_col20[1] <= data_out_4_20;
   result_col20[2] <= result_col20[1];
   result_col20[3] <= result_col20[2];
   result_col20[4] <= result_col20[3];
   result_col20[5] <= result_col20[4];
   result_col20[6] <= result_col20[5];
   result_col20[7] <= result_col20[6];
   result_col20[8] <= result_col20[7];
   result_col20[9] <= result_col20[8];
   result_col20[10] <= result_col20[9];
   result_col20[11] <= result_col20[10];
   result_col20[12] <= result_col20[11];
   result_col20[13] <= result_col20[12];
   result_col20[14] <= result_col20[13];
   result_col20[15] <= result_col20[14];
   result_col20[16] <= result_col20[15];
   result_col20[17] <= result_col20[16];
   result_col20[18] <= result_col20[17];
   result_col20[19] <= result_col20[18];
   result_col20[20] <= result_col20[19];
   result_col20[21] <= result_col20[20];
   result_col20[22] <= result_col20[21];
   result_col20[23] <= result_col20[22];
   result_col20[24] <= result_col20[23];
   result_col20[25] <= result_col20[24];
   result_col20[26] <= result_col20[25];
   result_col20[27] <= result_col20[26];
   result_col20[28] <= result_col20[27];
   result_col20[29] <= result_col20[28];
   result_col20[30] <= result_col20[29];
   result_col20[31] <= result_col20[30];
   result_col20[32] <= result_col20[31];
   result_col20[33] <= result_col20[32];
   result_col20[34] <= result_col20[33];
   result_col20[35] <= result_col20[34];
   result_col20[36] <= result_col20[35];
   result_col20[37] <= result_col20[36];
   result_col20[38] <= result_col20[37];
   result_col20[39] <= result_col20[38];
   result_col20[40] <= result_col20[39];
   result_col20[41] <= result_col20[40];
   result_col20[42] <= result_col20[41];
   result_col20[43] <= result_col20[42];
   result_col20[44] <= result_col20[43];
   result_col20[45] <= result_col20[44];
   result_col20[46] <= result_col20[45];
   result_col20[47] <= result_col20[46];
   result_col20[48] <= result_col20[47];
   result_col20[49] <= result_col20[48];
   result_col20[50] <= result_col20[49];
   result_col20[51] <= result_col20[50];
   result_col20[52] <= result_col20[51];
   result_col20[53] <= result_col20[52];
   result_col20[54] <= result_col20[53];
   result_col20[55] <= result_col20[54];
   result_col20[56] <= result_col20[55];
   result_col20[57] <= result_col20[56];
   result_col20[58] <= result_col20[57];
   result_col20[59] <= result_col20[58];
   result_col20[60] <= result_col20[59];
   result_col20[61] <= result_col20[60];
   result_col20[62] <= result_col20[61];
   result_col20[63] <= result_col20[62];
   result_col20[64] <= result_col20[63];
   result_col20[65] <= result_col20[64];
   result_col20[66] <= result_col20[65];
   result_col20[67] <= result_col20[66];
   result_col20[68] <= result_col20[67];
   result_col20[69] <= result_col20[68];
   result_col20[70] <= result_col20[69];
   result_col20[71] <= result_col20[70];
   result_col20[72] <= result_col20[71];
   result_col20[73] <= result_col20[72];
   result_col20[74] <= result_col20[73];
   result_col20[75] <= result_col20[74];
   result_col20[76] <= result_col20[75];
   result_col20[77] <= result_col20[76];
   result_col20[78] <= result_col20[77];
   result_col20[79] <= result_col20[78];
   result_col20[80] <= result_col20[79];
   result_col20[81] <= result_col20[80];
   result_col20[82] <= result_col20[81];
   result_col20[83] <= result_col20[82];
   result_col20[84] <= result_col20[83];
   result_col20[85] <= result_col20[84];
   result_col20[86] <= result_col20[85];
   result_col20[87] <= result_col20[86];
   result_col20[88] <= result_col20[87];
   result_col20[89] <= result_col20[88];
   result_col20[90] <= result_col20[89];
   result_col20[91] <= result_col20[90];
   result_col20[92] <= result_col20[91];
   result_col20[93] <= result_col20[92];
   result_col20[94] <= result_col20[93];
   result_col20[95] <= result_col20[94];
   result_col20[96] <= result_col20[95];
   result_col20[97] <= result_col20[96];
   result_col20[98] <= result_col20[97];
   result_col20[99] <= result_col20[98];
   result_col20[100] <= result_col20[99];
   result_col20[101] <= result_col20[100];
   result_col20[102] <= result_col20[101];
   result_col20[103] <= result_col20[102];
   result_col20[104] <= result_col20[103];
   result_col20[105] <= result_col20[104];
   result_col20[106] <= result_col20[105];
   result_col20[107] <= result_col20[106];
   result_col20[108] <= result_col20[107];
   result_col20[109] <= result_col20[108];
   result_col20[110] <= result_col20[109];
   result_col20[111] <= result_col20[110];
   result_col20[112] <= result_col20[111];
   result_col20[113] <= result_col20[112];
   result_col20[114] <= result_col20[113];
   result_col20[115] <= result_col20[114];
   result_col20[116] <= result_col20[115];
   result_col20[117] <= result_col20[116];
   result_col20[118] <= result_col20[117];
   result_col20[119] <= result_col20[118];
   result_col20[120] <= result_col20[119];
   result_col20[121] <= result_col20[120];
   result_col20[122] <= result_col20[121];
   result_col20[123] <= result_col20[122];
   result_col20[124] <= result_col20[123];
   result_col20[125] <= result_col20[124];
   result_col20[126] <= result_col20[125];
   result_col20[127] <= result_col20[126];
   result_col20[128] <= result_col20[127];
   result_col20[129] <= result_col20[128];
   result_col20[130] <= result_col20[129];
   result_col20[131] <= result_col20[130];
   result_col20[132] <= result_col20[131];
   result_col20[133] <= result_col20[132];
   result_col20[134] <= result_col20[133];
   result_col20[135] <= result_col20[134];
   result_col20[136] <= result_col20[135];
   result_col20[137] <= result_col20[136];
   result_col20[138] <= result_col20[137];
   result_col20[139] <= result_col20[138];
   result_col20[140] <= result_col20[139];
   result_col20[141] <= result_col20[140];
   result_col20[142] <= result_col20[141];
   result_col20[143] <= result_col20[142];
   result_col20[144] <= result_col20[143];
   result_col20[145] <= result_col20[144];
   result_col20[146] <= result_col20[145];

   result_col21[1] <= data_out_4_21;
   result_col21[2] <= result_col21[1];
   result_col21[3] <= result_col21[2];
   result_col21[4] <= result_col21[3];
   result_col21[5] <= result_col21[4];
   result_col21[6] <= result_col21[5];
   result_col21[7] <= result_col21[6];
   result_col21[8] <= result_col21[7];
   result_col21[9] <= result_col21[8];
   result_col21[10] <= result_col21[9];
   result_col21[11] <= result_col21[10];
   result_col21[12] <= result_col21[11];
   result_col21[13] <= result_col21[12];
   result_col21[14] <= result_col21[13];
   result_col21[15] <= result_col21[14];
   result_col21[16] <= result_col21[15];
   result_col21[17] <= result_col21[16];
   result_col21[18] <= result_col21[17];
   result_col21[19] <= result_col21[18];
   result_col21[20] <= result_col21[19];
   result_col21[21] <= result_col21[20];
   result_col21[22] <= result_col21[21];
   result_col21[23] <= result_col21[22];
   result_col21[24] <= result_col21[23];
   result_col21[25] <= result_col21[24];
   result_col21[26] <= result_col21[25];
   result_col21[27] <= result_col21[26];
   result_col21[28] <= result_col21[27];
   result_col21[29] <= result_col21[28];
   result_col21[30] <= result_col21[29];
   result_col21[31] <= result_col21[30];
   result_col21[32] <= result_col21[31];
   result_col21[33] <= result_col21[32];
   result_col21[34] <= result_col21[33];
   result_col21[35] <= result_col21[34];
   result_col21[36] <= result_col21[35];
   result_col21[37] <= result_col21[36];
   result_col21[38] <= result_col21[37];
   result_col21[39] <= result_col21[38];
   result_col21[40] <= result_col21[39];
   result_col21[41] <= result_col21[40];
   result_col21[42] <= result_col21[41];
   result_col21[43] <= result_col21[42];
   result_col21[44] <= result_col21[43];
   result_col21[45] <= result_col21[44];
   result_col21[46] <= result_col21[45];
   result_col21[47] <= result_col21[46];
   result_col21[48] <= result_col21[47];
   result_col21[49] <= result_col21[48];
   result_col21[50] <= result_col21[49];
   result_col21[51] <= result_col21[50];
   result_col21[52] <= result_col21[51];
   result_col21[53] <= result_col21[52];
   result_col21[54] <= result_col21[53];
   result_col21[55] <= result_col21[54];
   result_col21[56] <= result_col21[55];
   result_col21[57] <= result_col21[56];
   result_col21[58] <= result_col21[57];
   result_col21[59] <= result_col21[58];
   result_col21[60] <= result_col21[59];
   result_col21[61] <= result_col21[60];
   result_col21[62] <= result_col21[61];
   result_col21[63] <= result_col21[62];
   result_col21[64] <= result_col21[63];
   result_col21[65] <= result_col21[64];
   result_col21[66] <= result_col21[65];
   result_col21[67] <= result_col21[66];
   result_col21[68] <= result_col21[67];
   result_col21[69] <= result_col21[68];
   result_col21[70] <= result_col21[69];
   result_col21[71] <= result_col21[70];
   result_col21[72] <= result_col21[71];
   result_col21[73] <= result_col21[72];
   result_col21[74] <= result_col21[73];
   result_col21[75] <= result_col21[74];
   result_col21[76] <= result_col21[75];
   result_col21[77] <= result_col21[76];
   result_col21[78] <= result_col21[77];
   result_col21[79] <= result_col21[78];
   result_col21[80] <= result_col21[79];
   result_col21[81] <= result_col21[80];
   result_col21[82] <= result_col21[81];
   result_col21[83] <= result_col21[82];
   result_col21[84] <= result_col21[83];
   result_col21[85] <= result_col21[84];
   result_col21[86] <= result_col21[85];
   result_col21[87] <= result_col21[86];
   result_col21[88] <= result_col21[87];
   result_col21[89] <= result_col21[88];
   result_col21[90] <= result_col21[89];
   result_col21[91] <= result_col21[90];
   result_col21[92] <= result_col21[91];
   result_col21[93] <= result_col21[92];
   result_col21[94] <= result_col21[93];
   result_col21[95] <= result_col21[94];
   result_col21[96] <= result_col21[95];
   result_col21[97] <= result_col21[96];
   result_col21[98] <= result_col21[97];
   result_col21[99] <= result_col21[98];
   result_col21[100] <= result_col21[99];
   result_col21[101] <= result_col21[100];
   result_col21[102] <= result_col21[101];
   result_col21[103] <= result_col21[102];
   result_col21[104] <= result_col21[103];
   result_col21[105] <= result_col21[104];
   result_col21[106] <= result_col21[105];
   result_col21[107] <= result_col21[106];
   result_col21[108] <= result_col21[107];
   result_col21[109] <= result_col21[108];
   result_col21[110] <= result_col21[109];
   result_col21[111] <= result_col21[110];
   result_col21[112] <= result_col21[111];
   result_col21[113] <= result_col21[112];
   result_col21[114] <= result_col21[113];
   result_col21[115] <= result_col21[114];
   result_col21[116] <= result_col21[115];
   result_col21[117] <= result_col21[116];
   result_col21[118] <= result_col21[117];
   result_col21[119] <= result_col21[118];
   result_col21[120] <= result_col21[119];
   result_col21[121] <= result_col21[120];
   result_col21[122] <= result_col21[121];
   result_col21[123] <= result_col21[122];
   result_col21[124] <= result_col21[123];
   result_col21[125] <= result_col21[124];
   result_col21[126] <= result_col21[125];
   result_col21[127] <= result_col21[126];
   result_col21[128] <= result_col21[127];
   result_col21[129] <= result_col21[128];
   result_col21[130] <= result_col21[129];
   result_col21[131] <= result_col21[130];
   result_col21[132] <= result_col21[131];
   result_col21[133] <= result_col21[132];
   result_col21[134] <= result_col21[133];
   result_col21[135] <= result_col21[134];
   result_col21[136] <= result_col21[135];
   result_col21[137] <= result_col21[136];
   result_col21[138] <= result_col21[137];
   result_col21[139] <= result_col21[138];
   result_col21[140] <= result_col21[139];
   result_col21[141] <= result_col21[140];
   result_col21[142] <= result_col21[141];
   result_col21[143] <= result_col21[142];
   result_col21[144] <= result_col21[143];
   result_col21[145] <= result_col21[144];

   result_col22[1] <= data_out_4_22;
   result_col22[2] <= result_col22[1];
   result_col22[3] <= result_col22[2];
   result_col22[4] <= result_col22[3];
   result_col22[5] <= result_col22[4];
   result_col22[6] <= result_col22[5];
   result_col22[7] <= result_col22[6];
   result_col22[8] <= result_col22[7];
   result_col22[9] <= result_col22[8];
   result_col22[10] <= result_col22[9];
   result_col22[11] <= result_col22[10];
   result_col22[12] <= result_col22[11];
   result_col22[13] <= result_col22[12];
   result_col22[14] <= result_col22[13];
   result_col22[15] <= result_col22[14];
   result_col22[16] <= result_col22[15];
   result_col22[17] <= result_col22[16];
   result_col22[18] <= result_col22[17];
   result_col22[19] <= result_col22[18];
   result_col22[20] <= result_col22[19];
   result_col22[21] <= result_col22[20];
   result_col22[22] <= result_col22[21];
   result_col22[23] <= result_col22[22];
   result_col22[24] <= result_col22[23];
   result_col22[25] <= result_col22[24];
   result_col22[26] <= result_col22[25];
   result_col22[27] <= result_col22[26];
   result_col22[28] <= result_col22[27];
   result_col22[29] <= result_col22[28];
   result_col22[30] <= result_col22[29];
   result_col22[31] <= result_col22[30];
   result_col22[32] <= result_col22[31];
   result_col22[33] <= result_col22[32];
   result_col22[34] <= result_col22[33];
   result_col22[35] <= result_col22[34];
   result_col22[36] <= result_col22[35];
   result_col22[37] <= result_col22[36];
   result_col22[38] <= result_col22[37];
   result_col22[39] <= result_col22[38];
   result_col22[40] <= result_col22[39];
   result_col22[41] <= result_col22[40];
   result_col22[42] <= result_col22[41];
   result_col22[43] <= result_col22[42];
   result_col22[44] <= result_col22[43];
   result_col22[45] <= result_col22[44];
   result_col22[46] <= result_col22[45];
   result_col22[47] <= result_col22[46];
   result_col22[48] <= result_col22[47];
   result_col22[49] <= result_col22[48];
   result_col22[50] <= result_col22[49];
   result_col22[51] <= result_col22[50];
   result_col22[52] <= result_col22[51];
   result_col22[53] <= result_col22[52];
   result_col22[54] <= result_col22[53];
   result_col22[55] <= result_col22[54];
   result_col22[56] <= result_col22[55];
   result_col22[57] <= result_col22[56];
   result_col22[58] <= result_col22[57];
   result_col22[59] <= result_col22[58];
   result_col22[60] <= result_col22[59];
   result_col22[61] <= result_col22[60];
   result_col22[62] <= result_col22[61];
   result_col22[63] <= result_col22[62];
   result_col22[64] <= result_col22[63];
   result_col22[65] <= result_col22[64];
   result_col22[66] <= result_col22[65];
   result_col22[67] <= result_col22[66];
   result_col22[68] <= result_col22[67];
   result_col22[69] <= result_col22[68];
   result_col22[70] <= result_col22[69];
   result_col22[71] <= result_col22[70];
   result_col22[72] <= result_col22[71];
   result_col22[73] <= result_col22[72];
   result_col22[74] <= result_col22[73];
   result_col22[75] <= result_col22[74];
   result_col22[76] <= result_col22[75];
   result_col22[77] <= result_col22[76];
   result_col22[78] <= result_col22[77];
   result_col22[79] <= result_col22[78];
   result_col22[80] <= result_col22[79];
   result_col22[81] <= result_col22[80];
   result_col22[82] <= result_col22[81];
   result_col22[83] <= result_col22[82];
   result_col22[84] <= result_col22[83];
   result_col22[85] <= result_col22[84];
   result_col22[86] <= result_col22[85];
   result_col22[87] <= result_col22[86];
   result_col22[88] <= result_col22[87];
   result_col22[89] <= result_col22[88];
   result_col22[90] <= result_col22[89];
   result_col22[91] <= result_col22[90];
   result_col22[92] <= result_col22[91];
   result_col22[93] <= result_col22[92];
   result_col22[94] <= result_col22[93];
   result_col22[95] <= result_col22[94];
   result_col22[96] <= result_col22[95];
   result_col22[97] <= result_col22[96];
   result_col22[98] <= result_col22[97];
   result_col22[99] <= result_col22[98];
   result_col22[100] <= result_col22[99];
   result_col22[101] <= result_col22[100];
   result_col22[102] <= result_col22[101];
   result_col22[103] <= result_col22[102];
   result_col22[104] <= result_col22[103];
   result_col22[105] <= result_col22[104];
   result_col22[106] <= result_col22[105];
   result_col22[107] <= result_col22[106];
   result_col22[108] <= result_col22[107];
   result_col22[109] <= result_col22[108];
   result_col22[110] <= result_col22[109];
   result_col22[111] <= result_col22[110];
   result_col22[112] <= result_col22[111];
   result_col22[113] <= result_col22[112];
   result_col22[114] <= result_col22[113];
   result_col22[115] <= result_col22[114];
   result_col22[116] <= result_col22[115];
   result_col22[117] <= result_col22[116];
   result_col22[118] <= result_col22[117];
   result_col22[119] <= result_col22[118];
   result_col22[120] <= result_col22[119];
   result_col22[121] <= result_col22[120];
   result_col22[122] <= result_col22[121];
   result_col22[123] <= result_col22[122];
   result_col22[124] <= result_col22[123];
   result_col22[125] <= result_col22[124];
   result_col22[126] <= result_col22[125];
   result_col22[127] <= result_col22[126];
   result_col22[128] <= result_col22[127];
   result_col22[129] <= result_col22[128];
   result_col22[130] <= result_col22[129];
   result_col22[131] <= result_col22[130];
   result_col22[132] <= result_col22[131];
   result_col22[133] <= result_col22[132];
   result_col22[134] <= result_col22[133];
   result_col22[135] <= result_col22[134];
   result_col22[136] <= result_col22[135];
   result_col22[137] <= result_col22[136];
   result_col22[138] <= result_col22[137];
   result_col22[139] <= result_col22[138];
   result_col22[140] <= result_col22[139];
   result_col22[141] <= result_col22[140];
   result_col22[142] <= result_col22[141];
   result_col22[143] <= result_col22[142];
   result_col22[144] <= result_col22[143];

   result_col23[1] <= data_out_4_23;
   result_col23[2] <= result_col23[1];
   result_col23[3] <= result_col23[2];
   result_col23[4] <= result_col23[3];
   result_col23[5] <= result_col23[4];
   result_col23[6] <= result_col23[5];
   result_col23[7] <= result_col23[6];
   result_col23[8] <= result_col23[7];
   result_col23[9] <= result_col23[8];
   result_col23[10] <= result_col23[9];
   result_col23[11] <= result_col23[10];
   result_col23[12] <= result_col23[11];
   result_col23[13] <= result_col23[12];
   result_col23[14] <= result_col23[13];
   result_col23[15] <= result_col23[14];
   result_col23[16] <= result_col23[15];
   result_col23[17] <= result_col23[16];
   result_col23[18] <= result_col23[17];
   result_col23[19] <= result_col23[18];
   result_col23[20] <= result_col23[19];
   result_col23[21] <= result_col23[20];
   result_col23[22] <= result_col23[21];
   result_col23[23] <= result_col23[22];
   result_col23[24] <= result_col23[23];
   result_col23[25] <= result_col23[24];
   result_col23[26] <= result_col23[25];
   result_col23[27] <= result_col23[26];
   result_col23[28] <= result_col23[27];
   result_col23[29] <= result_col23[28];
   result_col23[30] <= result_col23[29];
   result_col23[31] <= result_col23[30];
   result_col23[32] <= result_col23[31];
   result_col23[33] <= result_col23[32];
   result_col23[34] <= result_col23[33];
   result_col23[35] <= result_col23[34];
   result_col23[36] <= result_col23[35];
   result_col23[37] <= result_col23[36];
   result_col23[38] <= result_col23[37];
   result_col23[39] <= result_col23[38];
   result_col23[40] <= result_col23[39];
   result_col23[41] <= result_col23[40];
   result_col23[42] <= result_col23[41];
   result_col23[43] <= result_col23[42];
   result_col23[44] <= result_col23[43];
   result_col23[45] <= result_col23[44];
   result_col23[46] <= result_col23[45];
   result_col23[47] <= result_col23[46];
   result_col23[48] <= result_col23[47];
   result_col23[49] <= result_col23[48];
   result_col23[50] <= result_col23[49];
   result_col23[51] <= result_col23[50];
   result_col23[52] <= result_col23[51];
   result_col23[53] <= result_col23[52];
   result_col23[54] <= result_col23[53];
   result_col23[55] <= result_col23[54];
   result_col23[56] <= result_col23[55];
   result_col23[57] <= result_col23[56];
   result_col23[58] <= result_col23[57];
   result_col23[59] <= result_col23[58];
   result_col23[60] <= result_col23[59];
   result_col23[61] <= result_col23[60];
   result_col23[62] <= result_col23[61];
   result_col23[63] <= result_col23[62];
   result_col23[64] <= result_col23[63];
   result_col23[65] <= result_col23[64];
   result_col23[66] <= result_col23[65];
   result_col23[67] <= result_col23[66];
   result_col23[68] <= result_col23[67];
   result_col23[69] <= result_col23[68];
   result_col23[70] <= result_col23[69];
   result_col23[71] <= result_col23[70];
   result_col23[72] <= result_col23[71];
   result_col23[73] <= result_col23[72];
   result_col23[74] <= result_col23[73];
   result_col23[75] <= result_col23[74];
   result_col23[76] <= result_col23[75];
   result_col23[77] <= result_col23[76];
   result_col23[78] <= result_col23[77];
   result_col23[79] <= result_col23[78];
   result_col23[80] <= result_col23[79];
   result_col23[81] <= result_col23[80];
   result_col23[82] <= result_col23[81];
   result_col23[83] <= result_col23[82];
   result_col23[84] <= result_col23[83];
   result_col23[85] <= result_col23[84];
   result_col23[86] <= result_col23[85];
   result_col23[87] <= result_col23[86];
   result_col23[88] <= result_col23[87];
   result_col23[89] <= result_col23[88];
   result_col23[90] <= result_col23[89];
   result_col23[91] <= result_col23[90];
   result_col23[92] <= result_col23[91];
   result_col23[93] <= result_col23[92];
   result_col23[94] <= result_col23[93];
   result_col23[95] <= result_col23[94];
   result_col23[96] <= result_col23[95];
   result_col23[97] <= result_col23[96];
   result_col23[98] <= result_col23[97];
   result_col23[99] <= result_col23[98];
   result_col23[100] <= result_col23[99];
   result_col23[101] <= result_col23[100];
   result_col23[102] <= result_col23[101];
   result_col23[103] <= result_col23[102];
   result_col23[104] <= result_col23[103];
   result_col23[105] <= result_col23[104];
   result_col23[106] <= result_col23[105];
   result_col23[107] <= result_col23[106];
   result_col23[108] <= result_col23[107];
   result_col23[109] <= result_col23[108];
   result_col23[110] <= result_col23[109];
   result_col23[111] <= result_col23[110];
   result_col23[112] <= result_col23[111];
   result_col23[113] <= result_col23[112];
   result_col23[114] <= result_col23[113];
   result_col23[115] <= result_col23[114];
   result_col23[116] <= result_col23[115];
   result_col23[117] <= result_col23[116];
   result_col23[118] <= result_col23[117];
   result_col23[119] <= result_col23[118];
   result_col23[120] <= result_col23[119];
   result_col23[121] <= result_col23[120];
   result_col23[122] <= result_col23[121];
   result_col23[123] <= result_col23[122];
   result_col23[124] <= result_col23[123];
   result_col23[125] <= result_col23[124];
   result_col23[126] <= result_col23[125];
   result_col23[127] <= result_col23[126];
   result_col23[128] <= result_col23[127];
   result_col23[129] <= result_col23[128];
   result_col23[130] <= result_col23[129];
   result_col23[131] <= result_col23[130];
   result_col23[132] <= result_col23[131];
   result_col23[133] <= result_col23[132];
   result_col23[134] <= result_col23[133];
   result_col23[135] <= result_col23[134];
   result_col23[136] <= result_col23[135];
   result_col23[137] <= result_col23[136];
   result_col23[138] <= result_col23[137];
   result_col23[139] <= result_col23[138];
   result_col23[140] <= result_col23[139];
   result_col23[141] <= result_col23[140];
   result_col23[142] <= result_col23[141];
   result_col23[143] <= result_col23[142];

   result_col24[1] <= data_out_4_24;
   result_col24[2] <= result_col24[1];
   result_col24[3] <= result_col24[2];
   result_col24[4] <= result_col24[3];
   result_col24[5] <= result_col24[4];
   result_col24[6] <= result_col24[5];
   result_col24[7] <= result_col24[6];
   result_col24[8] <= result_col24[7];
   result_col24[9] <= result_col24[8];
   result_col24[10] <= result_col24[9];
   result_col24[11] <= result_col24[10];
   result_col24[12] <= result_col24[11];
   result_col24[13] <= result_col24[12];
   result_col24[14] <= result_col24[13];
   result_col24[15] <= result_col24[14];
   result_col24[16] <= result_col24[15];
   result_col24[17] <= result_col24[16];
   result_col24[18] <= result_col24[17];
   result_col24[19] <= result_col24[18];
   result_col24[20] <= result_col24[19];
   result_col24[21] <= result_col24[20];
   result_col24[22] <= result_col24[21];
   result_col24[23] <= result_col24[22];
   result_col24[24] <= result_col24[23];
   result_col24[25] <= result_col24[24];
   result_col24[26] <= result_col24[25];
   result_col24[27] <= result_col24[26];
   result_col24[28] <= result_col24[27];
   result_col24[29] <= result_col24[28];
   result_col24[30] <= result_col24[29];
   result_col24[31] <= result_col24[30];
   result_col24[32] <= result_col24[31];
   result_col24[33] <= result_col24[32];
   result_col24[34] <= result_col24[33];
   result_col24[35] <= result_col24[34];
   result_col24[36] <= result_col24[35];
   result_col24[37] <= result_col24[36];
   result_col24[38] <= result_col24[37];
   result_col24[39] <= result_col24[38];
   result_col24[40] <= result_col24[39];
   result_col24[41] <= result_col24[40];
   result_col24[42] <= result_col24[41];
   result_col24[43] <= result_col24[42];
   result_col24[44] <= result_col24[43];
   result_col24[45] <= result_col24[44];
   result_col24[46] <= result_col24[45];
   result_col24[47] <= result_col24[46];
   result_col24[48] <= result_col24[47];
   result_col24[49] <= result_col24[48];
   result_col24[50] <= result_col24[49];
   result_col24[51] <= result_col24[50];
   result_col24[52] <= result_col24[51];
   result_col24[53] <= result_col24[52];
   result_col24[54] <= result_col24[53];
   result_col24[55] <= result_col24[54];
   result_col24[56] <= result_col24[55];
   result_col24[57] <= result_col24[56];
   result_col24[58] <= result_col24[57];
   result_col24[59] <= result_col24[58];
   result_col24[60] <= result_col24[59];
   result_col24[61] <= result_col24[60];
   result_col24[62] <= result_col24[61];
   result_col24[63] <= result_col24[62];
   result_col24[64] <= result_col24[63];
   result_col24[65] <= result_col24[64];
   result_col24[66] <= result_col24[65];
   result_col24[67] <= result_col24[66];
   result_col24[68] <= result_col24[67];
   result_col24[69] <= result_col24[68];
   result_col24[70] <= result_col24[69];
   result_col24[71] <= result_col24[70];
   result_col24[72] <= result_col24[71];
   result_col24[73] <= result_col24[72];
   result_col24[74] <= result_col24[73];
   result_col24[75] <= result_col24[74];
   result_col24[76] <= result_col24[75];
   result_col24[77] <= result_col24[76];
   result_col24[78] <= result_col24[77];
   result_col24[79] <= result_col24[78];
   result_col24[80] <= result_col24[79];
   result_col24[81] <= result_col24[80];
   result_col24[82] <= result_col24[81];
   result_col24[83] <= result_col24[82];
   result_col24[84] <= result_col24[83];
   result_col24[85] <= result_col24[84];
   result_col24[86] <= result_col24[85];
   result_col24[87] <= result_col24[86];
   result_col24[88] <= result_col24[87];
   result_col24[89] <= result_col24[88];
   result_col24[90] <= result_col24[89];
   result_col24[91] <= result_col24[90];
   result_col24[92] <= result_col24[91];
   result_col24[93] <= result_col24[92];
   result_col24[94] <= result_col24[93];
   result_col24[95] <= result_col24[94];
   result_col24[96] <= result_col24[95];
   result_col24[97] <= result_col24[96];
   result_col24[98] <= result_col24[97];
   result_col24[99] <= result_col24[98];
   result_col24[100] <= result_col24[99];
   result_col24[101] <= result_col24[100];
   result_col24[102] <= result_col24[101];
   result_col24[103] <= result_col24[102];
   result_col24[104] <= result_col24[103];
   result_col24[105] <= result_col24[104];
   result_col24[106] <= result_col24[105];
   result_col24[107] <= result_col24[106];
   result_col24[108] <= result_col24[107];
   result_col24[109] <= result_col24[108];
   result_col24[110] <= result_col24[109];
   result_col24[111] <= result_col24[110];
   result_col24[112] <= result_col24[111];
   result_col24[113] <= result_col24[112];
   result_col24[114] <= result_col24[113];
   result_col24[115] <= result_col24[114];
   result_col24[116] <= result_col24[115];
   result_col24[117] <= result_col24[116];
   result_col24[118] <= result_col24[117];
   result_col24[119] <= result_col24[118];
   result_col24[120] <= result_col24[119];
   result_col24[121] <= result_col24[120];
   result_col24[122] <= result_col24[121];
   result_col24[123] <= result_col24[122];
   result_col24[124] <= result_col24[123];
   result_col24[125] <= result_col24[124];
   result_col24[126] <= result_col24[125];
   result_col24[127] <= result_col24[126];
   result_col24[128] <= result_col24[127];
   result_col24[129] <= result_col24[128];
   result_col24[130] <= result_col24[129];
   result_col24[131] <= result_col24[130];
   result_col24[132] <= result_col24[131];
   result_col24[133] <= result_col24[132];
   result_col24[134] <= result_col24[133];
   result_col24[135] <= result_col24[134];
   result_col24[136] <= result_col24[135];
   result_col24[137] <= result_col24[136];
   result_col24[138] <= result_col24[137];
   result_col24[139] <= result_col24[138];
   result_col24[140] <= result_col24[139];
   result_col24[141] <= result_col24[140];
   result_col24[142] <= result_col24[141];

   result_col25[1] <= data_out_4_25;
   result_col25[2] <= result_col25[1];
   result_col25[3] <= result_col25[2];
   result_col25[4] <= result_col25[3];
   result_col25[5] <= result_col25[4];
   result_col25[6] <= result_col25[5];
   result_col25[7] <= result_col25[6];
   result_col25[8] <= result_col25[7];
   result_col25[9] <= result_col25[8];
   result_col25[10] <= result_col25[9];
   result_col25[11] <= result_col25[10];
   result_col25[12] <= result_col25[11];
   result_col25[13] <= result_col25[12];
   result_col25[14] <= result_col25[13];
   result_col25[15] <= result_col25[14];
   result_col25[16] <= result_col25[15];
   result_col25[17] <= result_col25[16];
   result_col25[18] <= result_col25[17];
   result_col25[19] <= result_col25[18];
   result_col25[20] <= result_col25[19];
   result_col25[21] <= result_col25[20];
   result_col25[22] <= result_col25[21];
   result_col25[23] <= result_col25[22];
   result_col25[24] <= result_col25[23];
   result_col25[25] <= result_col25[24];
   result_col25[26] <= result_col25[25];
   result_col25[27] <= result_col25[26];
   result_col25[28] <= result_col25[27];
   result_col25[29] <= result_col25[28];
   result_col25[30] <= result_col25[29];
   result_col25[31] <= result_col25[30];
   result_col25[32] <= result_col25[31];
   result_col25[33] <= result_col25[32];
   result_col25[34] <= result_col25[33];
   result_col25[35] <= result_col25[34];
   result_col25[36] <= result_col25[35];
   result_col25[37] <= result_col25[36];
   result_col25[38] <= result_col25[37];
   result_col25[39] <= result_col25[38];
   result_col25[40] <= result_col25[39];
   result_col25[41] <= result_col25[40];
   result_col25[42] <= result_col25[41];
   result_col25[43] <= result_col25[42];
   result_col25[44] <= result_col25[43];
   result_col25[45] <= result_col25[44];
   result_col25[46] <= result_col25[45];
   result_col25[47] <= result_col25[46];
   result_col25[48] <= result_col25[47];
   result_col25[49] <= result_col25[48];
   result_col25[50] <= result_col25[49];
   result_col25[51] <= result_col25[50];
   result_col25[52] <= result_col25[51];
   result_col25[53] <= result_col25[52];
   result_col25[54] <= result_col25[53];
   result_col25[55] <= result_col25[54];
   result_col25[56] <= result_col25[55];
   result_col25[57] <= result_col25[56];
   result_col25[58] <= result_col25[57];
   result_col25[59] <= result_col25[58];
   result_col25[60] <= result_col25[59];
   result_col25[61] <= result_col25[60];
   result_col25[62] <= result_col25[61];
   result_col25[63] <= result_col25[62];
   result_col25[64] <= result_col25[63];
   result_col25[65] <= result_col25[64];
   result_col25[66] <= result_col25[65];
   result_col25[67] <= result_col25[66];
   result_col25[68] <= result_col25[67];
   result_col25[69] <= result_col25[68];
   result_col25[70] <= result_col25[69];
   result_col25[71] <= result_col25[70];
   result_col25[72] <= result_col25[71];
   result_col25[73] <= result_col25[72];
   result_col25[74] <= result_col25[73];
   result_col25[75] <= result_col25[74];
   result_col25[76] <= result_col25[75];
   result_col25[77] <= result_col25[76];
   result_col25[78] <= result_col25[77];
   result_col25[79] <= result_col25[78];
   result_col25[80] <= result_col25[79];
   result_col25[81] <= result_col25[80];
   result_col25[82] <= result_col25[81];
   result_col25[83] <= result_col25[82];
   result_col25[84] <= result_col25[83];
   result_col25[85] <= result_col25[84];
   result_col25[86] <= result_col25[85];
   result_col25[87] <= result_col25[86];
   result_col25[88] <= result_col25[87];
   result_col25[89] <= result_col25[88];
   result_col25[90] <= result_col25[89];
   result_col25[91] <= result_col25[90];
   result_col25[92] <= result_col25[91];
   result_col25[93] <= result_col25[92];
   result_col25[94] <= result_col25[93];
   result_col25[95] <= result_col25[94];
   result_col25[96] <= result_col25[95];
   result_col25[97] <= result_col25[96];
   result_col25[98] <= result_col25[97];
   result_col25[99] <= result_col25[98];
   result_col25[100] <= result_col25[99];
   result_col25[101] <= result_col25[100];
   result_col25[102] <= result_col25[101];
   result_col25[103] <= result_col25[102];
   result_col25[104] <= result_col25[103];
   result_col25[105] <= result_col25[104];
   result_col25[106] <= result_col25[105];
   result_col25[107] <= result_col25[106];
   result_col25[108] <= result_col25[107];
   result_col25[109] <= result_col25[108];
   result_col25[110] <= result_col25[109];
   result_col25[111] <= result_col25[110];
   result_col25[112] <= result_col25[111];
   result_col25[113] <= result_col25[112];
   result_col25[114] <= result_col25[113];
   result_col25[115] <= result_col25[114];
   result_col25[116] <= result_col25[115];
   result_col25[117] <= result_col25[116];
   result_col25[118] <= result_col25[117];
   result_col25[119] <= result_col25[118];
   result_col25[120] <= result_col25[119];
   result_col25[121] <= result_col25[120];
   result_col25[122] <= result_col25[121];
   result_col25[123] <= result_col25[122];
   result_col25[124] <= result_col25[123];
   result_col25[125] <= result_col25[124];
   result_col25[126] <= result_col25[125];
   result_col25[127] <= result_col25[126];
   result_col25[128] <= result_col25[127];
   result_col25[129] <= result_col25[128];
   result_col25[130] <= result_col25[129];
   result_col25[131] <= result_col25[130];
   result_col25[132] <= result_col25[131];
   result_col25[133] <= result_col25[132];
   result_col25[134] <= result_col25[133];
   result_col25[135] <= result_col25[134];
   result_col25[136] <= result_col25[135];
   result_col25[137] <= result_col25[136];
   result_col25[138] <= result_col25[137];
   result_col25[139] <= result_col25[138];
   result_col25[140] <= result_col25[139];
   result_col25[141] <= result_col25[140];

   result_col26[1] <= data_out_4_26;
   result_col26[2] <= result_col26[1];
   result_col26[3] <= result_col26[2];
   result_col26[4] <= result_col26[3];
   result_col26[5] <= result_col26[4];
   result_col26[6] <= result_col26[5];
   result_col26[7] <= result_col26[6];
   result_col26[8] <= result_col26[7];
   result_col26[9] <= result_col26[8];
   result_col26[10] <= result_col26[9];
   result_col26[11] <= result_col26[10];
   result_col26[12] <= result_col26[11];
   result_col26[13] <= result_col26[12];
   result_col26[14] <= result_col26[13];
   result_col26[15] <= result_col26[14];
   result_col26[16] <= result_col26[15];
   result_col26[17] <= result_col26[16];
   result_col26[18] <= result_col26[17];
   result_col26[19] <= result_col26[18];
   result_col26[20] <= result_col26[19];
   result_col26[21] <= result_col26[20];
   result_col26[22] <= result_col26[21];
   result_col26[23] <= result_col26[22];
   result_col26[24] <= result_col26[23];
   result_col26[25] <= result_col26[24];
   result_col26[26] <= result_col26[25];
   result_col26[27] <= result_col26[26];
   result_col26[28] <= result_col26[27];
   result_col26[29] <= result_col26[28];
   result_col26[30] <= result_col26[29];
   result_col26[31] <= result_col26[30];
   result_col26[32] <= result_col26[31];
   result_col26[33] <= result_col26[32];
   result_col26[34] <= result_col26[33];
   result_col26[35] <= result_col26[34];
   result_col26[36] <= result_col26[35];
   result_col26[37] <= result_col26[36];
   result_col26[38] <= result_col26[37];
   result_col26[39] <= result_col26[38];
   result_col26[40] <= result_col26[39];
   result_col26[41] <= result_col26[40];
   result_col26[42] <= result_col26[41];
   result_col26[43] <= result_col26[42];
   result_col26[44] <= result_col26[43];
   result_col26[45] <= result_col26[44];
   result_col26[46] <= result_col26[45];
   result_col26[47] <= result_col26[46];
   result_col26[48] <= result_col26[47];
   result_col26[49] <= result_col26[48];
   result_col26[50] <= result_col26[49];
   result_col26[51] <= result_col26[50];
   result_col26[52] <= result_col26[51];
   result_col26[53] <= result_col26[52];
   result_col26[54] <= result_col26[53];
   result_col26[55] <= result_col26[54];
   result_col26[56] <= result_col26[55];
   result_col26[57] <= result_col26[56];
   result_col26[58] <= result_col26[57];
   result_col26[59] <= result_col26[58];
   result_col26[60] <= result_col26[59];
   result_col26[61] <= result_col26[60];
   result_col26[62] <= result_col26[61];
   result_col26[63] <= result_col26[62];
   result_col26[64] <= result_col26[63];
   result_col26[65] <= result_col26[64];
   result_col26[66] <= result_col26[65];
   result_col26[67] <= result_col26[66];
   result_col26[68] <= result_col26[67];
   result_col26[69] <= result_col26[68];
   result_col26[70] <= result_col26[69];
   result_col26[71] <= result_col26[70];
   result_col26[72] <= result_col26[71];
   result_col26[73] <= result_col26[72];
   result_col26[74] <= result_col26[73];
   result_col26[75] <= result_col26[74];
   result_col26[76] <= result_col26[75];
   result_col26[77] <= result_col26[76];
   result_col26[78] <= result_col26[77];
   result_col26[79] <= result_col26[78];
   result_col26[80] <= result_col26[79];
   result_col26[81] <= result_col26[80];
   result_col26[82] <= result_col26[81];
   result_col26[83] <= result_col26[82];
   result_col26[84] <= result_col26[83];
   result_col26[85] <= result_col26[84];
   result_col26[86] <= result_col26[85];
   result_col26[87] <= result_col26[86];
   result_col26[88] <= result_col26[87];
   result_col26[89] <= result_col26[88];
   result_col26[90] <= result_col26[89];
   result_col26[91] <= result_col26[90];
   result_col26[92] <= result_col26[91];
   result_col26[93] <= result_col26[92];
   result_col26[94] <= result_col26[93];
   result_col26[95] <= result_col26[94];
   result_col26[96] <= result_col26[95];
   result_col26[97] <= result_col26[96];
   result_col26[98] <= result_col26[97];
   result_col26[99] <= result_col26[98];
   result_col26[100] <= result_col26[99];
   result_col26[101] <= result_col26[100];
   result_col26[102] <= result_col26[101];
   result_col26[103] <= result_col26[102];
   result_col26[104] <= result_col26[103];
   result_col26[105] <= result_col26[104];
   result_col26[106] <= result_col26[105];
   result_col26[107] <= result_col26[106];
   result_col26[108] <= result_col26[107];
   result_col26[109] <= result_col26[108];
   result_col26[110] <= result_col26[109];
   result_col26[111] <= result_col26[110];
   result_col26[112] <= result_col26[111];
   result_col26[113] <= result_col26[112];
   result_col26[114] <= result_col26[113];
   result_col26[115] <= result_col26[114];
   result_col26[116] <= result_col26[115];
   result_col26[117] <= result_col26[116];
   result_col26[118] <= result_col26[117];
   result_col26[119] <= result_col26[118];
   result_col26[120] <= result_col26[119];
   result_col26[121] <= result_col26[120];
   result_col26[122] <= result_col26[121];
   result_col26[123] <= result_col26[122];
   result_col26[124] <= result_col26[123];
   result_col26[125] <= result_col26[124];
   result_col26[126] <= result_col26[125];
   result_col26[127] <= result_col26[126];
   result_col26[128] <= result_col26[127];
   result_col26[129] <= result_col26[128];
   result_col26[130] <= result_col26[129];
   result_col26[131] <= result_col26[130];
   result_col26[132] <= result_col26[131];
   result_col26[133] <= result_col26[132];
   result_col26[134] <= result_col26[133];
   result_col26[135] <= result_col26[134];
   result_col26[136] <= result_col26[135];
   result_col26[137] <= result_col26[136];
   result_col26[138] <= result_col26[137];
   result_col26[139] <= result_col26[138];
   result_col26[140] <= result_col26[139];

   result_col27[1] <= data_out_4_27;
   result_col27[2] <= result_col27[1];
   result_col27[3] <= result_col27[2];
   result_col27[4] <= result_col27[3];
   result_col27[5] <= result_col27[4];
   result_col27[6] <= result_col27[5];
   result_col27[7] <= result_col27[6];
   result_col27[8] <= result_col27[7];
   result_col27[9] <= result_col27[8];
   result_col27[10] <= result_col27[9];
   result_col27[11] <= result_col27[10];
   result_col27[12] <= result_col27[11];
   result_col27[13] <= result_col27[12];
   result_col27[14] <= result_col27[13];
   result_col27[15] <= result_col27[14];
   result_col27[16] <= result_col27[15];
   result_col27[17] <= result_col27[16];
   result_col27[18] <= result_col27[17];
   result_col27[19] <= result_col27[18];
   result_col27[20] <= result_col27[19];
   result_col27[21] <= result_col27[20];
   result_col27[22] <= result_col27[21];
   result_col27[23] <= result_col27[22];
   result_col27[24] <= result_col27[23];
   result_col27[25] <= result_col27[24];
   result_col27[26] <= result_col27[25];
   result_col27[27] <= result_col27[26];
   result_col27[28] <= result_col27[27];
   result_col27[29] <= result_col27[28];
   result_col27[30] <= result_col27[29];
   result_col27[31] <= result_col27[30];
   result_col27[32] <= result_col27[31];
   result_col27[33] <= result_col27[32];
   result_col27[34] <= result_col27[33];
   result_col27[35] <= result_col27[34];
   result_col27[36] <= result_col27[35];
   result_col27[37] <= result_col27[36];
   result_col27[38] <= result_col27[37];
   result_col27[39] <= result_col27[38];
   result_col27[40] <= result_col27[39];
   result_col27[41] <= result_col27[40];
   result_col27[42] <= result_col27[41];
   result_col27[43] <= result_col27[42];
   result_col27[44] <= result_col27[43];
   result_col27[45] <= result_col27[44];
   result_col27[46] <= result_col27[45];
   result_col27[47] <= result_col27[46];
   result_col27[48] <= result_col27[47];
   result_col27[49] <= result_col27[48];
   result_col27[50] <= result_col27[49];
   result_col27[51] <= result_col27[50];
   result_col27[52] <= result_col27[51];
   result_col27[53] <= result_col27[52];
   result_col27[54] <= result_col27[53];
   result_col27[55] <= result_col27[54];
   result_col27[56] <= result_col27[55];
   result_col27[57] <= result_col27[56];
   result_col27[58] <= result_col27[57];
   result_col27[59] <= result_col27[58];
   result_col27[60] <= result_col27[59];
   result_col27[61] <= result_col27[60];
   result_col27[62] <= result_col27[61];
   result_col27[63] <= result_col27[62];
   result_col27[64] <= result_col27[63];
   result_col27[65] <= result_col27[64];
   result_col27[66] <= result_col27[65];
   result_col27[67] <= result_col27[66];
   result_col27[68] <= result_col27[67];
   result_col27[69] <= result_col27[68];
   result_col27[70] <= result_col27[69];
   result_col27[71] <= result_col27[70];
   result_col27[72] <= result_col27[71];
   result_col27[73] <= result_col27[72];
   result_col27[74] <= result_col27[73];
   result_col27[75] <= result_col27[74];
   result_col27[76] <= result_col27[75];
   result_col27[77] <= result_col27[76];
   result_col27[78] <= result_col27[77];
   result_col27[79] <= result_col27[78];
   result_col27[80] <= result_col27[79];
   result_col27[81] <= result_col27[80];
   result_col27[82] <= result_col27[81];
   result_col27[83] <= result_col27[82];
   result_col27[84] <= result_col27[83];
   result_col27[85] <= result_col27[84];
   result_col27[86] <= result_col27[85];
   result_col27[87] <= result_col27[86];
   result_col27[88] <= result_col27[87];
   result_col27[89] <= result_col27[88];
   result_col27[90] <= result_col27[89];
   result_col27[91] <= result_col27[90];
   result_col27[92] <= result_col27[91];
   result_col27[93] <= result_col27[92];
   result_col27[94] <= result_col27[93];
   result_col27[95] <= result_col27[94];
   result_col27[96] <= result_col27[95];
   result_col27[97] <= result_col27[96];
   result_col27[98] <= result_col27[97];
   result_col27[99] <= result_col27[98];
   result_col27[100] <= result_col27[99];
   result_col27[101] <= result_col27[100];
   result_col27[102] <= result_col27[101];
   result_col27[103] <= result_col27[102];
   result_col27[104] <= result_col27[103];
   result_col27[105] <= result_col27[104];
   result_col27[106] <= result_col27[105];
   result_col27[107] <= result_col27[106];
   result_col27[108] <= result_col27[107];
   result_col27[109] <= result_col27[108];
   result_col27[110] <= result_col27[109];
   result_col27[111] <= result_col27[110];
   result_col27[112] <= result_col27[111];
   result_col27[113] <= result_col27[112];
   result_col27[114] <= result_col27[113];
   result_col27[115] <= result_col27[114];
   result_col27[116] <= result_col27[115];
   result_col27[117] <= result_col27[116];
   result_col27[118] <= result_col27[117];
   result_col27[119] <= result_col27[118];
   result_col27[120] <= result_col27[119];
   result_col27[121] <= result_col27[120];
   result_col27[122] <= result_col27[121];
   result_col27[123] <= result_col27[122];
   result_col27[124] <= result_col27[123];
   result_col27[125] <= result_col27[124];
   result_col27[126] <= result_col27[125];
   result_col27[127] <= result_col27[126];
   result_col27[128] <= result_col27[127];
   result_col27[129] <= result_col27[128];
   result_col27[130] <= result_col27[129];
   result_col27[131] <= result_col27[130];
   result_col27[132] <= result_col27[131];
   result_col27[133] <= result_col27[132];
   result_col27[134] <= result_col27[133];
   result_col27[135] <= result_col27[134];
   result_col27[136] <= result_col27[135];
   result_col27[137] <= result_col27[136];
   result_col27[138] <= result_col27[137];
   result_col27[139] <= result_col27[138];

   result_col28[1] <= data_out_4_28;
   result_col28[2] <= result_col28[1];
   result_col28[3] <= result_col28[2];
   result_col28[4] <= result_col28[3];
   result_col28[5] <= result_col28[4];
   result_col28[6] <= result_col28[5];
   result_col28[7] <= result_col28[6];
   result_col28[8] <= result_col28[7];
   result_col28[9] <= result_col28[8];
   result_col28[10] <= result_col28[9];
   result_col28[11] <= result_col28[10];
   result_col28[12] <= result_col28[11];
   result_col28[13] <= result_col28[12];
   result_col28[14] <= result_col28[13];
   result_col28[15] <= result_col28[14];
   result_col28[16] <= result_col28[15];
   result_col28[17] <= result_col28[16];
   result_col28[18] <= result_col28[17];
   result_col28[19] <= result_col28[18];
   result_col28[20] <= result_col28[19];
   result_col28[21] <= result_col28[20];
   result_col28[22] <= result_col28[21];
   result_col28[23] <= result_col28[22];
   result_col28[24] <= result_col28[23];
   result_col28[25] <= result_col28[24];
   result_col28[26] <= result_col28[25];
   result_col28[27] <= result_col28[26];
   result_col28[28] <= result_col28[27];
   result_col28[29] <= result_col28[28];
   result_col28[30] <= result_col28[29];
   result_col28[31] <= result_col28[30];
   result_col28[32] <= result_col28[31];
   result_col28[33] <= result_col28[32];
   result_col28[34] <= result_col28[33];
   result_col28[35] <= result_col28[34];
   result_col28[36] <= result_col28[35];
   result_col28[37] <= result_col28[36];
   result_col28[38] <= result_col28[37];
   result_col28[39] <= result_col28[38];
   result_col28[40] <= result_col28[39];
   result_col28[41] <= result_col28[40];
   result_col28[42] <= result_col28[41];
   result_col28[43] <= result_col28[42];
   result_col28[44] <= result_col28[43];
   result_col28[45] <= result_col28[44];
   result_col28[46] <= result_col28[45];
   result_col28[47] <= result_col28[46];
   result_col28[48] <= result_col28[47];
   result_col28[49] <= result_col28[48];
   result_col28[50] <= result_col28[49];
   result_col28[51] <= result_col28[50];
   result_col28[52] <= result_col28[51];
   result_col28[53] <= result_col28[52];
   result_col28[54] <= result_col28[53];
   result_col28[55] <= result_col28[54];
   result_col28[56] <= result_col28[55];
   result_col28[57] <= result_col28[56];
   result_col28[58] <= result_col28[57];
   result_col28[59] <= result_col28[58];
   result_col28[60] <= result_col28[59];
   result_col28[61] <= result_col28[60];
   result_col28[62] <= result_col28[61];
   result_col28[63] <= result_col28[62];
   result_col28[64] <= result_col28[63];
   result_col28[65] <= result_col28[64];
   result_col28[66] <= result_col28[65];
   result_col28[67] <= result_col28[66];
   result_col28[68] <= result_col28[67];
   result_col28[69] <= result_col28[68];
   result_col28[70] <= result_col28[69];
   result_col28[71] <= result_col28[70];
   result_col28[72] <= result_col28[71];
   result_col28[73] <= result_col28[72];
   result_col28[74] <= result_col28[73];
   result_col28[75] <= result_col28[74];
   result_col28[76] <= result_col28[75];
   result_col28[77] <= result_col28[76];
   result_col28[78] <= result_col28[77];
   result_col28[79] <= result_col28[78];
   result_col28[80] <= result_col28[79];
   result_col28[81] <= result_col28[80];
   result_col28[82] <= result_col28[81];
   result_col28[83] <= result_col28[82];
   result_col28[84] <= result_col28[83];
   result_col28[85] <= result_col28[84];
   result_col28[86] <= result_col28[85];
   result_col28[87] <= result_col28[86];
   result_col28[88] <= result_col28[87];
   result_col28[89] <= result_col28[88];
   result_col28[90] <= result_col28[89];
   result_col28[91] <= result_col28[90];
   result_col28[92] <= result_col28[91];
   result_col28[93] <= result_col28[92];
   result_col28[94] <= result_col28[93];
   result_col28[95] <= result_col28[94];
   result_col28[96] <= result_col28[95];
   result_col28[97] <= result_col28[96];
   result_col28[98] <= result_col28[97];
   result_col28[99] <= result_col28[98];
   result_col28[100] <= result_col28[99];
   result_col28[101] <= result_col28[100];
   result_col28[102] <= result_col28[101];
   result_col28[103] <= result_col28[102];
   result_col28[104] <= result_col28[103];
   result_col28[105] <= result_col28[104];
   result_col28[106] <= result_col28[105];
   result_col28[107] <= result_col28[106];
   result_col28[108] <= result_col28[107];
   result_col28[109] <= result_col28[108];
   result_col28[110] <= result_col28[109];
   result_col28[111] <= result_col28[110];
   result_col28[112] <= result_col28[111];
   result_col28[113] <= result_col28[112];
   result_col28[114] <= result_col28[113];
   result_col28[115] <= result_col28[114];
   result_col28[116] <= result_col28[115];
   result_col28[117] <= result_col28[116];
   result_col28[118] <= result_col28[117];
   result_col28[119] <= result_col28[118];
   result_col28[120] <= result_col28[119];
   result_col28[121] <= result_col28[120];
   result_col28[122] <= result_col28[121];
   result_col28[123] <= result_col28[122];
   result_col28[124] <= result_col28[123];
   result_col28[125] <= result_col28[124];
   result_col28[126] <= result_col28[125];
   result_col28[127] <= result_col28[126];
   result_col28[128] <= result_col28[127];
   result_col28[129] <= result_col28[128];
   result_col28[130] <= result_col28[129];
   result_col28[131] <= result_col28[130];
   result_col28[132] <= result_col28[131];
   result_col28[133] <= result_col28[132];
   result_col28[134] <= result_col28[133];
   result_col28[135] <= result_col28[134];
   result_col28[136] <= result_col28[135];
   result_col28[137] <= result_col28[136];
   result_col28[138] <= result_col28[137];

   result_col29[1] <= data_out_4_29;
   result_col29[2] <= result_col29[1];
   result_col29[3] <= result_col29[2];
   result_col29[4] <= result_col29[3];
   result_col29[5] <= result_col29[4];
   result_col29[6] <= result_col29[5];
   result_col29[7] <= result_col29[6];
   result_col29[8] <= result_col29[7];
   result_col29[9] <= result_col29[8];
   result_col29[10] <= result_col29[9];
   result_col29[11] <= result_col29[10];
   result_col29[12] <= result_col29[11];
   result_col29[13] <= result_col29[12];
   result_col29[14] <= result_col29[13];
   result_col29[15] <= result_col29[14];
   result_col29[16] <= result_col29[15];
   result_col29[17] <= result_col29[16];
   result_col29[18] <= result_col29[17];
   result_col29[19] <= result_col29[18];
   result_col29[20] <= result_col29[19];
   result_col29[21] <= result_col29[20];
   result_col29[22] <= result_col29[21];
   result_col29[23] <= result_col29[22];
   result_col29[24] <= result_col29[23];
   result_col29[25] <= result_col29[24];
   result_col29[26] <= result_col29[25];
   result_col29[27] <= result_col29[26];
   result_col29[28] <= result_col29[27];
   result_col29[29] <= result_col29[28];
   result_col29[30] <= result_col29[29];
   result_col29[31] <= result_col29[30];
   result_col29[32] <= result_col29[31];
   result_col29[33] <= result_col29[32];
   result_col29[34] <= result_col29[33];
   result_col29[35] <= result_col29[34];
   result_col29[36] <= result_col29[35];
   result_col29[37] <= result_col29[36];
   result_col29[38] <= result_col29[37];
   result_col29[39] <= result_col29[38];
   result_col29[40] <= result_col29[39];
   result_col29[41] <= result_col29[40];
   result_col29[42] <= result_col29[41];
   result_col29[43] <= result_col29[42];
   result_col29[44] <= result_col29[43];
   result_col29[45] <= result_col29[44];
   result_col29[46] <= result_col29[45];
   result_col29[47] <= result_col29[46];
   result_col29[48] <= result_col29[47];
   result_col29[49] <= result_col29[48];
   result_col29[50] <= result_col29[49];
   result_col29[51] <= result_col29[50];
   result_col29[52] <= result_col29[51];
   result_col29[53] <= result_col29[52];
   result_col29[54] <= result_col29[53];
   result_col29[55] <= result_col29[54];
   result_col29[56] <= result_col29[55];
   result_col29[57] <= result_col29[56];
   result_col29[58] <= result_col29[57];
   result_col29[59] <= result_col29[58];
   result_col29[60] <= result_col29[59];
   result_col29[61] <= result_col29[60];
   result_col29[62] <= result_col29[61];
   result_col29[63] <= result_col29[62];
   result_col29[64] <= result_col29[63];
   result_col29[65] <= result_col29[64];
   result_col29[66] <= result_col29[65];
   result_col29[67] <= result_col29[66];
   result_col29[68] <= result_col29[67];
   result_col29[69] <= result_col29[68];
   result_col29[70] <= result_col29[69];
   result_col29[71] <= result_col29[70];
   result_col29[72] <= result_col29[71];
   result_col29[73] <= result_col29[72];
   result_col29[74] <= result_col29[73];
   result_col29[75] <= result_col29[74];
   result_col29[76] <= result_col29[75];
   result_col29[77] <= result_col29[76];
   result_col29[78] <= result_col29[77];
   result_col29[79] <= result_col29[78];
   result_col29[80] <= result_col29[79];
   result_col29[81] <= result_col29[80];
   result_col29[82] <= result_col29[81];
   result_col29[83] <= result_col29[82];
   result_col29[84] <= result_col29[83];
   result_col29[85] <= result_col29[84];
   result_col29[86] <= result_col29[85];
   result_col29[87] <= result_col29[86];
   result_col29[88] <= result_col29[87];
   result_col29[89] <= result_col29[88];
   result_col29[90] <= result_col29[89];
   result_col29[91] <= result_col29[90];
   result_col29[92] <= result_col29[91];
   result_col29[93] <= result_col29[92];
   result_col29[94] <= result_col29[93];
   result_col29[95] <= result_col29[94];
   result_col29[96] <= result_col29[95];
   result_col29[97] <= result_col29[96];
   result_col29[98] <= result_col29[97];
   result_col29[99] <= result_col29[98];
   result_col29[100] <= result_col29[99];
   result_col29[101] <= result_col29[100];
   result_col29[102] <= result_col29[101];
   result_col29[103] <= result_col29[102];
   result_col29[104] <= result_col29[103];
   result_col29[105] <= result_col29[104];
   result_col29[106] <= result_col29[105];
   result_col29[107] <= result_col29[106];
   result_col29[108] <= result_col29[107];
   result_col29[109] <= result_col29[108];
   result_col29[110] <= result_col29[109];
   result_col29[111] <= result_col29[110];
   result_col29[112] <= result_col29[111];
   result_col29[113] <= result_col29[112];
   result_col29[114] <= result_col29[113];
   result_col29[115] <= result_col29[114];
   result_col29[116] <= result_col29[115];
   result_col29[117] <= result_col29[116];
   result_col29[118] <= result_col29[117];
   result_col29[119] <= result_col29[118];
   result_col29[120] <= result_col29[119];
   result_col29[121] <= result_col29[120];
   result_col29[122] <= result_col29[121];
   result_col29[123] <= result_col29[122];
   result_col29[124] <= result_col29[123];
   result_col29[125] <= result_col29[124];
   result_col29[126] <= result_col29[125];
   result_col29[127] <= result_col29[126];
   result_col29[128] <= result_col29[127];
   result_col29[129] <= result_col29[128];
   result_col29[130] <= result_col29[129];
   result_col29[131] <= result_col29[130];
   result_col29[132] <= result_col29[131];
   result_col29[133] <= result_col29[132];
   result_col29[134] <= result_col29[133];
   result_col29[135] <= result_col29[134];
   result_col29[136] <= result_col29[135];
   result_col29[137] <= result_col29[136];

   result_col30[1] <= data_out_4_30;
   result_col30[2] <= result_col30[1];
   result_col30[3] <= result_col30[2];
   result_col30[4] <= result_col30[3];
   result_col30[5] <= result_col30[4];
   result_col30[6] <= result_col30[5];
   result_col30[7] <= result_col30[6];
   result_col30[8] <= result_col30[7];
   result_col30[9] <= result_col30[8];
   result_col30[10] <= result_col30[9];
   result_col30[11] <= result_col30[10];
   result_col30[12] <= result_col30[11];
   result_col30[13] <= result_col30[12];
   result_col30[14] <= result_col30[13];
   result_col30[15] <= result_col30[14];
   result_col30[16] <= result_col30[15];
   result_col30[17] <= result_col30[16];
   result_col30[18] <= result_col30[17];
   result_col30[19] <= result_col30[18];
   result_col30[20] <= result_col30[19];
   result_col30[21] <= result_col30[20];
   result_col30[22] <= result_col30[21];
   result_col30[23] <= result_col30[22];
   result_col30[24] <= result_col30[23];
   result_col30[25] <= result_col30[24];
   result_col30[26] <= result_col30[25];
   result_col30[27] <= result_col30[26];
   result_col30[28] <= result_col30[27];
   result_col30[29] <= result_col30[28];
   result_col30[30] <= result_col30[29];
   result_col30[31] <= result_col30[30];
   result_col30[32] <= result_col30[31];
   result_col30[33] <= result_col30[32];
   result_col30[34] <= result_col30[33];
   result_col30[35] <= result_col30[34];
   result_col30[36] <= result_col30[35];
   result_col30[37] <= result_col30[36];
   result_col30[38] <= result_col30[37];
   result_col30[39] <= result_col30[38];
   result_col30[40] <= result_col30[39];
   result_col30[41] <= result_col30[40];
   result_col30[42] <= result_col30[41];
   result_col30[43] <= result_col30[42];
   result_col30[44] <= result_col30[43];
   result_col30[45] <= result_col30[44];
   result_col30[46] <= result_col30[45];
   result_col30[47] <= result_col30[46];
   result_col30[48] <= result_col30[47];
   result_col30[49] <= result_col30[48];
   result_col30[50] <= result_col30[49];
   result_col30[51] <= result_col30[50];
   result_col30[52] <= result_col30[51];
   result_col30[53] <= result_col30[52];
   result_col30[54] <= result_col30[53];
   result_col30[55] <= result_col30[54];
   result_col30[56] <= result_col30[55];
   result_col30[57] <= result_col30[56];
   result_col30[58] <= result_col30[57];
   result_col30[59] <= result_col30[58];
   result_col30[60] <= result_col30[59];
   result_col30[61] <= result_col30[60];
   result_col30[62] <= result_col30[61];
   result_col30[63] <= result_col30[62];
   result_col30[64] <= result_col30[63];
   result_col30[65] <= result_col30[64];
   result_col30[66] <= result_col30[65];
   result_col30[67] <= result_col30[66];
   result_col30[68] <= result_col30[67];
   result_col30[69] <= result_col30[68];
   result_col30[70] <= result_col30[69];
   result_col30[71] <= result_col30[70];
   result_col30[72] <= result_col30[71];
   result_col30[73] <= result_col30[72];
   result_col30[74] <= result_col30[73];
   result_col30[75] <= result_col30[74];
   result_col30[76] <= result_col30[75];
   result_col30[77] <= result_col30[76];
   result_col30[78] <= result_col30[77];
   result_col30[79] <= result_col30[78];
   result_col30[80] <= result_col30[79];
   result_col30[81] <= result_col30[80];
   result_col30[82] <= result_col30[81];
   result_col30[83] <= result_col30[82];
   result_col30[84] <= result_col30[83];
   result_col30[85] <= result_col30[84];
   result_col30[86] <= result_col30[85];
   result_col30[87] <= result_col30[86];
   result_col30[88] <= result_col30[87];
   result_col30[89] <= result_col30[88];
   result_col30[90] <= result_col30[89];
   result_col30[91] <= result_col30[90];
   result_col30[92] <= result_col30[91];
   result_col30[93] <= result_col30[92];
   result_col30[94] <= result_col30[93];
   result_col30[95] <= result_col30[94];
   result_col30[96] <= result_col30[95];
   result_col30[97] <= result_col30[96];
   result_col30[98] <= result_col30[97];
   result_col30[99] <= result_col30[98];
   result_col30[100] <= result_col30[99];
   result_col30[101] <= result_col30[100];
   result_col30[102] <= result_col30[101];
   result_col30[103] <= result_col30[102];
   result_col30[104] <= result_col30[103];
   result_col30[105] <= result_col30[104];
   result_col30[106] <= result_col30[105];
   result_col30[107] <= result_col30[106];
   result_col30[108] <= result_col30[107];
   result_col30[109] <= result_col30[108];
   result_col30[110] <= result_col30[109];
   result_col30[111] <= result_col30[110];
   result_col30[112] <= result_col30[111];
   result_col30[113] <= result_col30[112];
   result_col30[114] <= result_col30[113];
   result_col30[115] <= result_col30[114];
   result_col30[116] <= result_col30[115];
   result_col30[117] <= result_col30[116];
   result_col30[118] <= result_col30[117];
   result_col30[119] <= result_col30[118];
   result_col30[120] <= result_col30[119];
   result_col30[121] <= result_col30[120];
   result_col30[122] <= result_col30[121];
   result_col30[123] <= result_col30[122];
   result_col30[124] <= result_col30[123];
   result_col30[125] <= result_col30[124];
   result_col30[126] <= result_col30[125];
   result_col30[127] <= result_col30[126];
   result_col30[128] <= result_col30[127];
   result_col30[129] <= result_col30[128];
   result_col30[130] <= result_col30[129];
   result_col30[131] <= result_col30[130];
   result_col30[132] <= result_col30[131];
   result_col30[133] <= result_col30[132];
   result_col30[134] <= result_col30[133];
   result_col30[135] <= result_col30[134];
   result_col30[136] <= result_col30[135];

   result_col31[1] <= data_out_4_31;
   result_col31[2] <= result_col31[1];
   result_col31[3] <= result_col31[2];
   result_col31[4] <= result_col31[3];
   result_col31[5] <= result_col31[4];
   result_col31[6] <= result_col31[5];
   result_col31[7] <= result_col31[6];
   result_col31[8] <= result_col31[7];
   result_col31[9] <= result_col31[8];
   result_col31[10] <= result_col31[9];
   result_col31[11] <= result_col31[10];
   result_col31[12] <= result_col31[11];
   result_col31[13] <= result_col31[12];
   result_col31[14] <= result_col31[13];
   result_col31[15] <= result_col31[14];
   result_col31[16] <= result_col31[15];
   result_col31[17] <= result_col31[16];
   result_col31[18] <= result_col31[17];
   result_col31[19] <= result_col31[18];
   result_col31[20] <= result_col31[19];
   result_col31[21] <= result_col31[20];
   result_col31[22] <= result_col31[21];
   result_col31[23] <= result_col31[22];
   result_col31[24] <= result_col31[23];
   result_col31[25] <= result_col31[24];
   result_col31[26] <= result_col31[25];
   result_col31[27] <= result_col31[26];
   result_col31[28] <= result_col31[27];
   result_col31[29] <= result_col31[28];
   result_col31[30] <= result_col31[29];
   result_col31[31] <= result_col31[30];
   result_col31[32] <= result_col31[31];
   result_col31[33] <= result_col31[32];
   result_col31[34] <= result_col31[33];
   result_col31[35] <= result_col31[34];
   result_col31[36] <= result_col31[35];
   result_col31[37] <= result_col31[36];
   result_col31[38] <= result_col31[37];
   result_col31[39] <= result_col31[38];
   result_col31[40] <= result_col31[39];
   result_col31[41] <= result_col31[40];
   result_col31[42] <= result_col31[41];
   result_col31[43] <= result_col31[42];
   result_col31[44] <= result_col31[43];
   result_col31[45] <= result_col31[44];
   result_col31[46] <= result_col31[45];
   result_col31[47] <= result_col31[46];
   result_col31[48] <= result_col31[47];
   result_col31[49] <= result_col31[48];
   result_col31[50] <= result_col31[49];
   result_col31[51] <= result_col31[50];
   result_col31[52] <= result_col31[51];
   result_col31[53] <= result_col31[52];
   result_col31[54] <= result_col31[53];
   result_col31[55] <= result_col31[54];
   result_col31[56] <= result_col31[55];
   result_col31[57] <= result_col31[56];
   result_col31[58] <= result_col31[57];
   result_col31[59] <= result_col31[58];
   result_col31[60] <= result_col31[59];
   result_col31[61] <= result_col31[60];
   result_col31[62] <= result_col31[61];
   result_col31[63] <= result_col31[62];
   result_col31[64] <= result_col31[63];
   result_col31[65] <= result_col31[64];
   result_col31[66] <= result_col31[65];
   result_col31[67] <= result_col31[66];
   result_col31[68] <= result_col31[67];
   result_col31[69] <= result_col31[68];
   result_col31[70] <= result_col31[69];
   result_col31[71] <= result_col31[70];
   result_col31[72] <= result_col31[71];
   result_col31[73] <= result_col31[72];
   result_col31[74] <= result_col31[73];
   result_col31[75] <= result_col31[74];
   result_col31[76] <= result_col31[75];
   result_col31[77] <= result_col31[76];
   result_col31[78] <= result_col31[77];
   result_col31[79] <= result_col31[78];
   result_col31[80] <= result_col31[79];
   result_col31[81] <= result_col31[80];
   result_col31[82] <= result_col31[81];
   result_col31[83] <= result_col31[82];
   result_col31[84] <= result_col31[83];
   result_col31[85] <= result_col31[84];
   result_col31[86] <= result_col31[85];
   result_col31[87] <= result_col31[86];
   result_col31[88] <= result_col31[87];
   result_col31[89] <= result_col31[88];
   result_col31[90] <= result_col31[89];
   result_col31[91] <= result_col31[90];
   result_col31[92] <= result_col31[91];
   result_col31[93] <= result_col31[92];
   result_col31[94] <= result_col31[93];
   result_col31[95] <= result_col31[94];
   result_col31[96] <= result_col31[95];
   result_col31[97] <= result_col31[96];
   result_col31[98] <= result_col31[97];
   result_col31[99] <= result_col31[98];
   result_col31[100] <= result_col31[99];
   result_col31[101] <= result_col31[100];
   result_col31[102] <= result_col31[101];
   result_col31[103] <= result_col31[102];
   result_col31[104] <= result_col31[103];
   result_col31[105] <= result_col31[104];
   result_col31[106] <= result_col31[105];
   result_col31[107] <= result_col31[106];
   result_col31[108] <= result_col31[107];
   result_col31[109] <= result_col31[108];
   result_col31[110] <= result_col31[109];
   result_col31[111] <= result_col31[110];
   result_col31[112] <= result_col31[111];
   result_col31[113] <= result_col31[112];
   result_col31[114] <= result_col31[113];
   result_col31[115] <= result_col31[114];
   result_col31[116] <= result_col31[115];
   result_col31[117] <= result_col31[116];
   result_col31[118] <= result_col31[117];
   result_col31[119] <= result_col31[118];
   result_col31[120] <= result_col31[119];
   result_col31[121] <= result_col31[120];
   result_col31[122] <= result_col31[121];
   result_col31[123] <= result_col31[122];
   result_col31[124] <= result_col31[123];
   result_col31[125] <= result_col31[124];
   result_col31[126] <= result_col31[125];
   result_col31[127] <= result_col31[126];
   result_col31[128] <= result_col31[127];
   result_col31[129] <= result_col31[128];
   result_col31[130] <= result_col31[129];
   result_col31[131] <= result_col31[130];
   result_col31[132] <= result_col31[131];
   result_col31[133] <= result_col31[132];
   result_col31[134] <= result_col31[133];
   result_col31[135] <= result_col31[134];

   result_col32[1] <= data_out_4_32;
   result_col32[2] <= result_col32[1];
   result_col32[3] <= result_col32[2];
   result_col32[4] <= result_col32[3];
   result_col32[5] <= result_col32[4];
   result_col32[6] <= result_col32[5];
   result_col32[7] <= result_col32[6];
   result_col32[8] <= result_col32[7];
   result_col32[9] <= result_col32[8];
   result_col32[10] <= result_col32[9];
   result_col32[11] <= result_col32[10];
   result_col32[12] <= result_col32[11];
   result_col32[13] <= result_col32[12];
   result_col32[14] <= result_col32[13];
   result_col32[15] <= result_col32[14];
   result_col32[16] <= result_col32[15];
   result_col32[17] <= result_col32[16];
   result_col32[18] <= result_col32[17];
   result_col32[19] <= result_col32[18];
   result_col32[20] <= result_col32[19];
   result_col32[21] <= result_col32[20];
   result_col32[22] <= result_col32[21];
   result_col32[23] <= result_col32[22];
   result_col32[24] <= result_col32[23];
   result_col32[25] <= result_col32[24];
   result_col32[26] <= result_col32[25];
   result_col32[27] <= result_col32[26];
   result_col32[28] <= result_col32[27];
   result_col32[29] <= result_col32[28];
   result_col32[30] <= result_col32[29];
   result_col32[31] <= result_col32[30];
   result_col32[32] <= result_col32[31];
   result_col32[33] <= result_col32[32];
   result_col32[34] <= result_col32[33];
   result_col32[35] <= result_col32[34];
   result_col32[36] <= result_col32[35];
   result_col32[37] <= result_col32[36];
   result_col32[38] <= result_col32[37];
   result_col32[39] <= result_col32[38];
   result_col32[40] <= result_col32[39];
   result_col32[41] <= result_col32[40];
   result_col32[42] <= result_col32[41];
   result_col32[43] <= result_col32[42];
   result_col32[44] <= result_col32[43];
   result_col32[45] <= result_col32[44];
   result_col32[46] <= result_col32[45];
   result_col32[47] <= result_col32[46];
   result_col32[48] <= result_col32[47];
   result_col32[49] <= result_col32[48];
   result_col32[50] <= result_col32[49];
   result_col32[51] <= result_col32[50];
   result_col32[52] <= result_col32[51];
   result_col32[53] <= result_col32[52];
   result_col32[54] <= result_col32[53];
   result_col32[55] <= result_col32[54];
   result_col32[56] <= result_col32[55];
   result_col32[57] <= result_col32[56];
   result_col32[58] <= result_col32[57];
   result_col32[59] <= result_col32[58];
   result_col32[60] <= result_col32[59];
   result_col32[61] <= result_col32[60];
   result_col32[62] <= result_col32[61];
   result_col32[63] <= result_col32[62];
   result_col32[64] <= result_col32[63];
   result_col32[65] <= result_col32[64];
   result_col32[66] <= result_col32[65];
   result_col32[67] <= result_col32[66];
   result_col32[68] <= result_col32[67];
   result_col32[69] <= result_col32[68];
   result_col32[70] <= result_col32[69];
   result_col32[71] <= result_col32[70];
   result_col32[72] <= result_col32[71];
   result_col32[73] <= result_col32[72];
   result_col32[74] <= result_col32[73];
   result_col32[75] <= result_col32[74];
   result_col32[76] <= result_col32[75];
   result_col32[77] <= result_col32[76];
   result_col32[78] <= result_col32[77];
   result_col32[79] <= result_col32[78];
   result_col32[80] <= result_col32[79];
   result_col32[81] <= result_col32[80];
   result_col32[82] <= result_col32[81];
   result_col32[83] <= result_col32[82];
   result_col32[84] <= result_col32[83];
   result_col32[85] <= result_col32[84];
   result_col32[86] <= result_col32[85];
   result_col32[87] <= result_col32[86];
   result_col32[88] <= result_col32[87];
   result_col32[89] <= result_col32[88];
   result_col32[90] <= result_col32[89];
   result_col32[91] <= result_col32[90];
   result_col32[92] <= result_col32[91];
   result_col32[93] <= result_col32[92];
   result_col32[94] <= result_col32[93];
   result_col32[95] <= result_col32[94];
   result_col32[96] <= result_col32[95];
   result_col32[97] <= result_col32[96];
   result_col32[98] <= result_col32[97];
   result_col32[99] <= result_col32[98];
   result_col32[100] <= result_col32[99];
   result_col32[101] <= result_col32[100];
   result_col32[102] <= result_col32[101];
   result_col32[103] <= result_col32[102];
   result_col32[104] <= result_col32[103];
   result_col32[105] <= result_col32[104];
   result_col32[106] <= result_col32[105];
   result_col32[107] <= result_col32[106];
   result_col32[108] <= result_col32[107];
   result_col32[109] <= result_col32[108];
   result_col32[110] <= result_col32[109];
   result_col32[111] <= result_col32[110];
   result_col32[112] <= result_col32[111];
   result_col32[113] <= result_col32[112];
   result_col32[114] <= result_col32[113];
   result_col32[115] <= result_col32[114];
   result_col32[116] <= result_col32[115];
   result_col32[117] <= result_col32[116];
   result_col32[118] <= result_col32[117];
   result_col32[119] <= result_col32[118];
   result_col32[120] <= result_col32[119];
   result_col32[121] <= result_col32[120];
   result_col32[122] <= result_col32[121];
   result_col32[123] <= result_col32[122];
   result_col32[124] <= result_col32[123];
   result_col32[125] <= result_col32[124];
   result_col32[126] <= result_col32[125];
   result_col32[127] <= result_col32[126];
   result_col32[128] <= result_col32[127];
   result_col32[129] <= result_col32[128];
   result_col32[130] <= result_col32[129];
   result_col32[131] <= result_col32[130];
   result_col32[132] <= result_col32[131];
   result_col32[133] <= result_col32[132];
   result_col32[134] <= result_col32[133];

   result_col33[1] <= data_out_4_33;
   result_col33[2] <= result_col33[1];
   result_col33[3] <= result_col33[2];
   result_col33[4] <= result_col33[3];
   result_col33[5] <= result_col33[4];
   result_col33[6] <= result_col33[5];
   result_col33[7] <= result_col33[6];
   result_col33[8] <= result_col33[7];
   result_col33[9] <= result_col33[8];
   result_col33[10] <= result_col33[9];
   result_col33[11] <= result_col33[10];
   result_col33[12] <= result_col33[11];
   result_col33[13] <= result_col33[12];
   result_col33[14] <= result_col33[13];
   result_col33[15] <= result_col33[14];
   result_col33[16] <= result_col33[15];
   result_col33[17] <= result_col33[16];
   result_col33[18] <= result_col33[17];
   result_col33[19] <= result_col33[18];
   result_col33[20] <= result_col33[19];
   result_col33[21] <= result_col33[20];
   result_col33[22] <= result_col33[21];
   result_col33[23] <= result_col33[22];
   result_col33[24] <= result_col33[23];
   result_col33[25] <= result_col33[24];
   result_col33[26] <= result_col33[25];
   result_col33[27] <= result_col33[26];
   result_col33[28] <= result_col33[27];
   result_col33[29] <= result_col33[28];
   result_col33[30] <= result_col33[29];
   result_col33[31] <= result_col33[30];
   result_col33[32] <= result_col33[31];
   result_col33[33] <= result_col33[32];
   result_col33[34] <= result_col33[33];
   result_col33[35] <= result_col33[34];
   result_col33[36] <= result_col33[35];
   result_col33[37] <= result_col33[36];
   result_col33[38] <= result_col33[37];
   result_col33[39] <= result_col33[38];
   result_col33[40] <= result_col33[39];
   result_col33[41] <= result_col33[40];
   result_col33[42] <= result_col33[41];
   result_col33[43] <= result_col33[42];
   result_col33[44] <= result_col33[43];
   result_col33[45] <= result_col33[44];
   result_col33[46] <= result_col33[45];
   result_col33[47] <= result_col33[46];
   result_col33[48] <= result_col33[47];
   result_col33[49] <= result_col33[48];
   result_col33[50] <= result_col33[49];
   result_col33[51] <= result_col33[50];
   result_col33[52] <= result_col33[51];
   result_col33[53] <= result_col33[52];
   result_col33[54] <= result_col33[53];
   result_col33[55] <= result_col33[54];
   result_col33[56] <= result_col33[55];
   result_col33[57] <= result_col33[56];
   result_col33[58] <= result_col33[57];
   result_col33[59] <= result_col33[58];
   result_col33[60] <= result_col33[59];
   result_col33[61] <= result_col33[60];
   result_col33[62] <= result_col33[61];
   result_col33[63] <= result_col33[62];
   result_col33[64] <= result_col33[63];
   result_col33[65] <= result_col33[64];
   result_col33[66] <= result_col33[65];
   result_col33[67] <= result_col33[66];
   result_col33[68] <= result_col33[67];
   result_col33[69] <= result_col33[68];
   result_col33[70] <= result_col33[69];
   result_col33[71] <= result_col33[70];
   result_col33[72] <= result_col33[71];
   result_col33[73] <= result_col33[72];
   result_col33[74] <= result_col33[73];
   result_col33[75] <= result_col33[74];
   result_col33[76] <= result_col33[75];
   result_col33[77] <= result_col33[76];
   result_col33[78] <= result_col33[77];
   result_col33[79] <= result_col33[78];
   result_col33[80] <= result_col33[79];
   result_col33[81] <= result_col33[80];
   result_col33[82] <= result_col33[81];
   result_col33[83] <= result_col33[82];
   result_col33[84] <= result_col33[83];
   result_col33[85] <= result_col33[84];
   result_col33[86] <= result_col33[85];
   result_col33[87] <= result_col33[86];
   result_col33[88] <= result_col33[87];
   result_col33[89] <= result_col33[88];
   result_col33[90] <= result_col33[89];
   result_col33[91] <= result_col33[90];
   result_col33[92] <= result_col33[91];
   result_col33[93] <= result_col33[92];
   result_col33[94] <= result_col33[93];
   result_col33[95] <= result_col33[94];
   result_col33[96] <= result_col33[95];
   result_col33[97] <= result_col33[96];
   result_col33[98] <= result_col33[97];
   result_col33[99] <= result_col33[98];
   result_col33[100] <= result_col33[99];
   result_col33[101] <= result_col33[100];
   result_col33[102] <= result_col33[101];
   result_col33[103] <= result_col33[102];
   result_col33[104] <= result_col33[103];
   result_col33[105] <= result_col33[104];
   result_col33[106] <= result_col33[105];
   result_col33[107] <= result_col33[106];
   result_col33[108] <= result_col33[107];
   result_col33[109] <= result_col33[108];
   result_col33[110] <= result_col33[109];
   result_col33[111] <= result_col33[110];
   result_col33[112] <= result_col33[111];
   result_col33[113] <= result_col33[112];
   result_col33[114] <= result_col33[113];
   result_col33[115] <= result_col33[114];
   result_col33[116] <= result_col33[115];
   result_col33[117] <= result_col33[116];
   result_col33[118] <= result_col33[117];
   result_col33[119] <= result_col33[118];
   result_col33[120] <= result_col33[119];
   result_col33[121] <= result_col33[120];
   result_col33[122] <= result_col33[121];
   result_col33[123] <= result_col33[122];
   result_col33[124] <= result_col33[123];
   result_col33[125] <= result_col33[124];
   result_col33[126] <= result_col33[125];
   result_col33[127] <= result_col33[126];
   result_col33[128] <= result_col33[127];
   result_col33[129] <= result_col33[128];
   result_col33[130] <= result_col33[129];
   result_col33[131] <= result_col33[130];
   result_col33[132] <= result_col33[131];
   result_col33[133] <= result_col33[132];

   result_col34[1] <= data_out_4_34;
   result_col34[2] <= result_col34[1];
   result_col34[3] <= result_col34[2];
   result_col34[4] <= result_col34[3];
   result_col34[5] <= result_col34[4];
   result_col34[6] <= result_col34[5];
   result_col34[7] <= result_col34[6];
   result_col34[8] <= result_col34[7];
   result_col34[9] <= result_col34[8];
   result_col34[10] <= result_col34[9];
   result_col34[11] <= result_col34[10];
   result_col34[12] <= result_col34[11];
   result_col34[13] <= result_col34[12];
   result_col34[14] <= result_col34[13];
   result_col34[15] <= result_col34[14];
   result_col34[16] <= result_col34[15];
   result_col34[17] <= result_col34[16];
   result_col34[18] <= result_col34[17];
   result_col34[19] <= result_col34[18];
   result_col34[20] <= result_col34[19];
   result_col34[21] <= result_col34[20];
   result_col34[22] <= result_col34[21];
   result_col34[23] <= result_col34[22];
   result_col34[24] <= result_col34[23];
   result_col34[25] <= result_col34[24];
   result_col34[26] <= result_col34[25];
   result_col34[27] <= result_col34[26];
   result_col34[28] <= result_col34[27];
   result_col34[29] <= result_col34[28];
   result_col34[30] <= result_col34[29];
   result_col34[31] <= result_col34[30];
   result_col34[32] <= result_col34[31];
   result_col34[33] <= result_col34[32];
   result_col34[34] <= result_col34[33];
   result_col34[35] <= result_col34[34];
   result_col34[36] <= result_col34[35];
   result_col34[37] <= result_col34[36];
   result_col34[38] <= result_col34[37];
   result_col34[39] <= result_col34[38];
   result_col34[40] <= result_col34[39];
   result_col34[41] <= result_col34[40];
   result_col34[42] <= result_col34[41];
   result_col34[43] <= result_col34[42];
   result_col34[44] <= result_col34[43];
   result_col34[45] <= result_col34[44];
   result_col34[46] <= result_col34[45];
   result_col34[47] <= result_col34[46];
   result_col34[48] <= result_col34[47];
   result_col34[49] <= result_col34[48];
   result_col34[50] <= result_col34[49];
   result_col34[51] <= result_col34[50];
   result_col34[52] <= result_col34[51];
   result_col34[53] <= result_col34[52];
   result_col34[54] <= result_col34[53];
   result_col34[55] <= result_col34[54];
   result_col34[56] <= result_col34[55];
   result_col34[57] <= result_col34[56];
   result_col34[58] <= result_col34[57];
   result_col34[59] <= result_col34[58];
   result_col34[60] <= result_col34[59];
   result_col34[61] <= result_col34[60];
   result_col34[62] <= result_col34[61];
   result_col34[63] <= result_col34[62];
   result_col34[64] <= result_col34[63];
   result_col34[65] <= result_col34[64];
   result_col34[66] <= result_col34[65];
   result_col34[67] <= result_col34[66];
   result_col34[68] <= result_col34[67];
   result_col34[69] <= result_col34[68];
   result_col34[70] <= result_col34[69];
   result_col34[71] <= result_col34[70];
   result_col34[72] <= result_col34[71];
   result_col34[73] <= result_col34[72];
   result_col34[74] <= result_col34[73];
   result_col34[75] <= result_col34[74];
   result_col34[76] <= result_col34[75];
   result_col34[77] <= result_col34[76];
   result_col34[78] <= result_col34[77];
   result_col34[79] <= result_col34[78];
   result_col34[80] <= result_col34[79];
   result_col34[81] <= result_col34[80];
   result_col34[82] <= result_col34[81];
   result_col34[83] <= result_col34[82];
   result_col34[84] <= result_col34[83];
   result_col34[85] <= result_col34[84];
   result_col34[86] <= result_col34[85];
   result_col34[87] <= result_col34[86];
   result_col34[88] <= result_col34[87];
   result_col34[89] <= result_col34[88];
   result_col34[90] <= result_col34[89];
   result_col34[91] <= result_col34[90];
   result_col34[92] <= result_col34[91];
   result_col34[93] <= result_col34[92];
   result_col34[94] <= result_col34[93];
   result_col34[95] <= result_col34[94];
   result_col34[96] <= result_col34[95];
   result_col34[97] <= result_col34[96];
   result_col34[98] <= result_col34[97];
   result_col34[99] <= result_col34[98];
   result_col34[100] <= result_col34[99];
   result_col34[101] <= result_col34[100];
   result_col34[102] <= result_col34[101];
   result_col34[103] <= result_col34[102];
   result_col34[104] <= result_col34[103];
   result_col34[105] <= result_col34[104];
   result_col34[106] <= result_col34[105];
   result_col34[107] <= result_col34[106];
   result_col34[108] <= result_col34[107];
   result_col34[109] <= result_col34[108];
   result_col34[110] <= result_col34[109];
   result_col34[111] <= result_col34[110];
   result_col34[112] <= result_col34[111];
   result_col34[113] <= result_col34[112];
   result_col34[114] <= result_col34[113];
   result_col34[115] <= result_col34[114];
   result_col34[116] <= result_col34[115];
   result_col34[117] <= result_col34[116];
   result_col34[118] <= result_col34[117];
   result_col34[119] <= result_col34[118];
   result_col34[120] <= result_col34[119];
   result_col34[121] <= result_col34[120];
   result_col34[122] <= result_col34[121];
   result_col34[123] <= result_col34[122];
   result_col34[124] <= result_col34[123];
   result_col34[125] <= result_col34[124];
   result_col34[126] <= result_col34[125];
   result_col34[127] <= result_col34[126];
   result_col34[128] <= result_col34[127];
   result_col34[129] <= result_col34[128];
   result_col34[130] <= result_col34[129];
   result_col34[131] <= result_col34[130];
   result_col34[132] <= result_col34[131];

   result_col35[1] <= data_out_4_35;
   result_col35[2] <= result_col35[1];
   result_col35[3] <= result_col35[2];
   result_col35[4] <= result_col35[3];
   result_col35[5] <= result_col35[4];
   result_col35[6] <= result_col35[5];
   result_col35[7] <= result_col35[6];
   result_col35[8] <= result_col35[7];
   result_col35[9] <= result_col35[8];
   result_col35[10] <= result_col35[9];
   result_col35[11] <= result_col35[10];
   result_col35[12] <= result_col35[11];
   result_col35[13] <= result_col35[12];
   result_col35[14] <= result_col35[13];
   result_col35[15] <= result_col35[14];
   result_col35[16] <= result_col35[15];
   result_col35[17] <= result_col35[16];
   result_col35[18] <= result_col35[17];
   result_col35[19] <= result_col35[18];
   result_col35[20] <= result_col35[19];
   result_col35[21] <= result_col35[20];
   result_col35[22] <= result_col35[21];
   result_col35[23] <= result_col35[22];
   result_col35[24] <= result_col35[23];
   result_col35[25] <= result_col35[24];
   result_col35[26] <= result_col35[25];
   result_col35[27] <= result_col35[26];
   result_col35[28] <= result_col35[27];
   result_col35[29] <= result_col35[28];
   result_col35[30] <= result_col35[29];
   result_col35[31] <= result_col35[30];
   result_col35[32] <= result_col35[31];
   result_col35[33] <= result_col35[32];
   result_col35[34] <= result_col35[33];
   result_col35[35] <= result_col35[34];
   result_col35[36] <= result_col35[35];
   result_col35[37] <= result_col35[36];
   result_col35[38] <= result_col35[37];
   result_col35[39] <= result_col35[38];
   result_col35[40] <= result_col35[39];
   result_col35[41] <= result_col35[40];
   result_col35[42] <= result_col35[41];
   result_col35[43] <= result_col35[42];
   result_col35[44] <= result_col35[43];
   result_col35[45] <= result_col35[44];
   result_col35[46] <= result_col35[45];
   result_col35[47] <= result_col35[46];
   result_col35[48] <= result_col35[47];
   result_col35[49] <= result_col35[48];
   result_col35[50] <= result_col35[49];
   result_col35[51] <= result_col35[50];
   result_col35[52] <= result_col35[51];
   result_col35[53] <= result_col35[52];
   result_col35[54] <= result_col35[53];
   result_col35[55] <= result_col35[54];
   result_col35[56] <= result_col35[55];
   result_col35[57] <= result_col35[56];
   result_col35[58] <= result_col35[57];
   result_col35[59] <= result_col35[58];
   result_col35[60] <= result_col35[59];
   result_col35[61] <= result_col35[60];
   result_col35[62] <= result_col35[61];
   result_col35[63] <= result_col35[62];
   result_col35[64] <= result_col35[63];
   result_col35[65] <= result_col35[64];
   result_col35[66] <= result_col35[65];
   result_col35[67] <= result_col35[66];
   result_col35[68] <= result_col35[67];
   result_col35[69] <= result_col35[68];
   result_col35[70] <= result_col35[69];
   result_col35[71] <= result_col35[70];
   result_col35[72] <= result_col35[71];
   result_col35[73] <= result_col35[72];
   result_col35[74] <= result_col35[73];
   result_col35[75] <= result_col35[74];
   result_col35[76] <= result_col35[75];
   result_col35[77] <= result_col35[76];
   result_col35[78] <= result_col35[77];
   result_col35[79] <= result_col35[78];
   result_col35[80] <= result_col35[79];
   result_col35[81] <= result_col35[80];
   result_col35[82] <= result_col35[81];
   result_col35[83] <= result_col35[82];
   result_col35[84] <= result_col35[83];
   result_col35[85] <= result_col35[84];
   result_col35[86] <= result_col35[85];
   result_col35[87] <= result_col35[86];
   result_col35[88] <= result_col35[87];
   result_col35[89] <= result_col35[88];
   result_col35[90] <= result_col35[89];
   result_col35[91] <= result_col35[90];
   result_col35[92] <= result_col35[91];
   result_col35[93] <= result_col35[92];
   result_col35[94] <= result_col35[93];
   result_col35[95] <= result_col35[94];
   result_col35[96] <= result_col35[95];
   result_col35[97] <= result_col35[96];
   result_col35[98] <= result_col35[97];
   result_col35[99] <= result_col35[98];
   result_col35[100] <= result_col35[99];
   result_col35[101] <= result_col35[100];
   result_col35[102] <= result_col35[101];
   result_col35[103] <= result_col35[102];
   result_col35[104] <= result_col35[103];
   result_col35[105] <= result_col35[104];
   result_col35[106] <= result_col35[105];
   result_col35[107] <= result_col35[106];
   result_col35[108] <= result_col35[107];
   result_col35[109] <= result_col35[108];
   result_col35[110] <= result_col35[109];
   result_col35[111] <= result_col35[110];
   result_col35[112] <= result_col35[111];
   result_col35[113] <= result_col35[112];
   result_col35[114] <= result_col35[113];
   result_col35[115] <= result_col35[114];
   result_col35[116] <= result_col35[115];
   result_col35[117] <= result_col35[116];
   result_col35[118] <= result_col35[117];
   result_col35[119] <= result_col35[118];
   result_col35[120] <= result_col35[119];
   result_col35[121] <= result_col35[120];
   result_col35[122] <= result_col35[121];
   result_col35[123] <= result_col35[122];
   result_col35[124] <= result_col35[123];
   result_col35[125] <= result_col35[124];
   result_col35[126] <= result_col35[125];
   result_col35[127] <= result_col35[126];
   result_col35[128] <= result_col35[127];
   result_col35[129] <= result_col35[128];
   result_col35[130] <= result_col35[129];
   result_col35[131] <= result_col35[130];

   result_col36[1] <= data_out_4_36;
   result_col36[2] <= result_col36[1];
   result_col36[3] <= result_col36[2];
   result_col36[4] <= result_col36[3];
   result_col36[5] <= result_col36[4];
   result_col36[6] <= result_col36[5];
   result_col36[7] <= result_col36[6];
   result_col36[8] <= result_col36[7];
   result_col36[9] <= result_col36[8];
   result_col36[10] <= result_col36[9];
   result_col36[11] <= result_col36[10];
   result_col36[12] <= result_col36[11];
   result_col36[13] <= result_col36[12];
   result_col36[14] <= result_col36[13];
   result_col36[15] <= result_col36[14];
   result_col36[16] <= result_col36[15];
   result_col36[17] <= result_col36[16];
   result_col36[18] <= result_col36[17];
   result_col36[19] <= result_col36[18];
   result_col36[20] <= result_col36[19];
   result_col36[21] <= result_col36[20];
   result_col36[22] <= result_col36[21];
   result_col36[23] <= result_col36[22];
   result_col36[24] <= result_col36[23];
   result_col36[25] <= result_col36[24];
   result_col36[26] <= result_col36[25];
   result_col36[27] <= result_col36[26];
   result_col36[28] <= result_col36[27];
   result_col36[29] <= result_col36[28];
   result_col36[30] <= result_col36[29];
   result_col36[31] <= result_col36[30];
   result_col36[32] <= result_col36[31];
   result_col36[33] <= result_col36[32];
   result_col36[34] <= result_col36[33];
   result_col36[35] <= result_col36[34];
   result_col36[36] <= result_col36[35];
   result_col36[37] <= result_col36[36];
   result_col36[38] <= result_col36[37];
   result_col36[39] <= result_col36[38];
   result_col36[40] <= result_col36[39];
   result_col36[41] <= result_col36[40];
   result_col36[42] <= result_col36[41];
   result_col36[43] <= result_col36[42];
   result_col36[44] <= result_col36[43];
   result_col36[45] <= result_col36[44];
   result_col36[46] <= result_col36[45];
   result_col36[47] <= result_col36[46];
   result_col36[48] <= result_col36[47];
   result_col36[49] <= result_col36[48];
   result_col36[50] <= result_col36[49];
   result_col36[51] <= result_col36[50];
   result_col36[52] <= result_col36[51];
   result_col36[53] <= result_col36[52];
   result_col36[54] <= result_col36[53];
   result_col36[55] <= result_col36[54];
   result_col36[56] <= result_col36[55];
   result_col36[57] <= result_col36[56];
   result_col36[58] <= result_col36[57];
   result_col36[59] <= result_col36[58];
   result_col36[60] <= result_col36[59];
   result_col36[61] <= result_col36[60];
   result_col36[62] <= result_col36[61];
   result_col36[63] <= result_col36[62];
   result_col36[64] <= result_col36[63];
   result_col36[65] <= result_col36[64];
   result_col36[66] <= result_col36[65];
   result_col36[67] <= result_col36[66];
   result_col36[68] <= result_col36[67];
   result_col36[69] <= result_col36[68];
   result_col36[70] <= result_col36[69];
   result_col36[71] <= result_col36[70];
   result_col36[72] <= result_col36[71];
   result_col36[73] <= result_col36[72];
   result_col36[74] <= result_col36[73];
   result_col36[75] <= result_col36[74];
   result_col36[76] <= result_col36[75];
   result_col36[77] <= result_col36[76];
   result_col36[78] <= result_col36[77];
   result_col36[79] <= result_col36[78];
   result_col36[80] <= result_col36[79];
   result_col36[81] <= result_col36[80];
   result_col36[82] <= result_col36[81];
   result_col36[83] <= result_col36[82];
   result_col36[84] <= result_col36[83];
   result_col36[85] <= result_col36[84];
   result_col36[86] <= result_col36[85];
   result_col36[87] <= result_col36[86];
   result_col36[88] <= result_col36[87];
   result_col36[89] <= result_col36[88];
   result_col36[90] <= result_col36[89];
   result_col36[91] <= result_col36[90];
   result_col36[92] <= result_col36[91];
   result_col36[93] <= result_col36[92];
   result_col36[94] <= result_col36[93];
   result_col36[95] <= result_col36[94];
   result_col36[96] <= result_col36[95];
   result_col36[97] <= result_col36[96];
   result_col36[98] <= result_col36[97];
   result_col36[99] <= result_col36[98];
   result_col36[100] <= result_col36[99];
   result_col36[101] <= result_col36[100];
   result_col36[102] <= result_col36[101];
   result_col36[103] <= result_col36[102];
   result_col36[104] <= result_col36[103];
   result_col36[105] <= result_col36[104];
   result_col36[106] <= result_col36[105];
   result_col36[107] <= result_col36[106];
   result_col36[108] <= result_col36[107];
   result_col36[109] <= result_col36[108];
   result_col36[110] <= result_col36[109];
   result_col36[111] <= result_col36[110];
   result_col36[112] <= result_col36[111];
   result_col36[113] <= result_col36[112];
   result_col36[114] <= result_col36[113];
   result_col36[115] <= result_col36[114];
   result_col36[116] <= result_col36[115];
   result_col36[117] <= result_col36[116];
   result_col36[118] <= result_col36[117];
   result_col36[119] <= result_col36[118];
   result_col36[120] <= result_col36[119];
   result_col36[121] <= result_col36[120];
   result_col36[122] <= result_col36[121];
   result_col36[123] <= result_col36[122];
   result_col36[124] <= result_col36[123];
   result_col36[125] <= result_col36[124];
   result_col36[126] <= result_col36[125];
   result_col36[127] <= result_col36[126];
   result_col36[128] <= result_col36[127];
   result_col36[129] <= result_col36[128];
   result_col36[130] <= result_col36[129];

   result_col37[1] <= data_out_4_37;
   result_col37[2] <= result_col37[1];
   result_col37[3] <= result_col37[2];
   result_col37[4] <= result_col37[3];
   result_col37[5] <= result_col37[4];
   result_col37[6] <= result_col37[5];
   result_col37[7] <= result_col37[6];
   result_col37[8] <= result_col37[7];
   result_col37[9] <= result_col37[8];
   result_col37[10] <= result_col37[9];
   result_col37[11] <= result_col37[10];
   result_col37[12] <= result_col37[11];
   result_col37[13] <= result_col37[12];
   result_col37[14] <= result_col37[13];
   result_col37[15] <= result_col37[14];
   result_col37[16] <= result_col37[15];
   result_col37[17] <= result_col37[16];
   result_col37[18] <= result_col37[17];
   result_col37[19] <= result_col37[18];
   result_col37[20] <= result_col37[19];
   result_col37[21] <= result_col37[20];
   result_col37[22] <= result_col37[21];
   result_col37[23] <= result_col37[22];
   result_col37[24] <= result_col37[23];
   result_col37[25] <= result_col37[24];
   result_col37[26] <= result_col37[25];
   result_col37[27] <= result_col37[26];
   result_col37[28] <= result_col37[27];
   result_col37[29] <= result_col37[28];
   result_col37[30] <= result_col37[29];
   result_col37[31] <= result_col37[30];
   result_col37[32] <= result_col37[31];
   result_col37[33] <= result_col37[32];
   result_col37[34] <= result_col37[33];
   result_col37[35] <= result_col37[34];
   result_col37[36] <= result_col37[35];
   result_col37[37] <= result_col37[36];
   result_col37[38] <= result_col37[37];
   result_col37[39] <= result_col37[38];
   result_col37[40] <= result_col37[39];
   result_col37[41] <= result_col37[40];
   result_col37[42] <= result_col37[41];
   result_col37[43] <= result_col37[42];
   result_col37[44] <= result_col37[43];
   result_col37[45] <= result_col37[44];
   result_col37[46] <= result_col37[45];
   result_col37[47] <= result_col37[46];
   result_col37[48] <= result_col37[47];
   result_col37[49] <= result_col37[48];
   result_col37[50] <= result_col37[49];
   result_col37[51] <= result_col37[50];
   result_col37[52] <= result_col37[51];
   result_col37[53] <= result_col37[52];
   result_col37[54] <= result_col37[53];
   result_col37[55] <= result_col37[54];
   result_col37[56] <= result_col37[55];
   result_col37[57] <= result_col37[56];
   result_col37[58] <= result_col37[57];
   result_col37[59] <= result_col37[58];
   result_col37[60] <= result_col37[59];
   result_col37[61] <= result_col37[60];
   result_col37[62] <= result_col37[61];
   result_col37[63] <= result_col37[62];
   result_col37[64] <= result_col37[63];
   result_col37[65] <= result_col37[64];
   result_col37[66] <= result_col37[65];
   result_col37[67] <= result_col37[66];
   result_col37[68] <= result_col37[67];
   result_col37[69] <= result_col37[68];
   result_col37[70] <= result_col37[69];
   result_col37[71] <= result_col37[70];
   result_col37[72] <= result_col37[71];
   result_col37[73] <= result_col37[72];
   result_col37[74] <= result_col37[73];
   result_col37[75] <= result_col37[74];
   result_col37[76] <= result_col37[75];
   result_col37[77] <= result_col37[76];
   result_col37[78] <= result_col37[77];
   result_col37[79] <= result_col37[78];
   result_col37[80] <= result_col37[79];
   result_col37[81] <= result_col37[80];
   result_col37[82] <= result_col37[81];
   result_col37[83] <= result_col37[82];
   result_col37[84] <= result_col37[83];
   result_col37[85] <= result_col37[84];
   result_col37[86] <= result_col37[85];
   result_col37[87] <= result_col37[86];
   result_col37[88] <= result_col37[87];
   result_col37[89] <= result_col37[88];
   result_col37[90] <= result_col37[89];
   result_col37[91] <= result_col37[90];
   result_col37[92] <= result_col37[91];
   result_col37[93] <= result_col37[92];
   result_col37[94] <= result_col37[93];
   result_col37[95] <= result_col37[94];
   result_col37[96] <= result_col37[95];
   result_col37[97] <= result_col37[96];
   result_col37[98] <= result_col37[97];
   result_col37[99] <= result_col37[98];
   result_col37[100] <= result_col37[99];
   result_col37[101] <= result_col37[100];
   result_col37[102] <= result_col37[101];
   result_col37[103] <= result_col37[102];
   result_col37[104] <= result_col37[103];
   result_col37[105] <= result_col37[104];
   result_col37[106] <= result_col37[105];
   result_col37[107] <= result_col37[106];
   result_col37[108] <= result_col37[107];
   result_col37[109] <= result_col37[108];
   result_col37[110] <= result_col37[109];
   result_col37[111] <= result_col37[110];
   result_col37[112] <= result_col37[111];
   result_col37[113] <= result_col37[112];
   result_col37[114] <= result_col37[113];
   result_col37[115] <= result_col37[114];
   result_col37[116] <= result_col37[115];
   result_col37[117] <= result_col37[116];
   result_col37[118] <= result_col37[117];
   result_col37[119] <= result_col37[118];
   result_col37[120] <= result_col37[119];
   result_col37[121] <= result_col37[120];
   result_col37[122] <= result_col37[121];
   result_col37[123] <= result_col37[122];
   result_col37[124] <= result_col37[123];
   result_col37[125] <= result_col37[124];
   result_col37[126] <= result_col37[125];
   result_col37[127] <= result_col37[126];
   result_col37[128] <= result_col37[127];
   result_col37[129] <= result_col37[128];

   result_col38[1] <= data_out_4_38;
   result_col38[2] <= result_col38[1];
   result_col38[3] <= result_col38[2];
   result_col38[4] <= result_col38[3];
   result_col38[5] <= result_col38[4];
   result_col38[6] <= result_col38[5];
   result_col38[7] <= result_col38[6];
   result_col38[8] <= result_col38[7];
   result_col38[9] <= result_col38[8];
   result_col38[10] <= result_col38[9];
   result_col38[11] <= result_col38[10];
   result_col38[12] <= result_col38[11];
   result_col38[13] <= result_col38[12];
   result_col38[14] <= result_col38[13];
   result_col38[15] <= result_col38[14];
   result_col38[16] <= result_col38[15];
   result_col38[17] <= result_col38[16];
   result_col38[18] <= result_col38[17];
   result_col38[19] <= result_col38[18];
   result_col38[20] <= result_col38[19];
   result_col38[21] <= result_col38[20];
   result_col38[22] <= result_col38[21];
   result_col38[23] <= result_col38[22];
   result_col38[24] <= result_col38[23];
   result_col38[25] <= result_col38[24];
   result_col38[26] <= result_col38[25];
   result_col38[27] <= result_col38[26];
   result_col38[28] <= result_col38[27];
   result_col38[29] <= result_col38[28];
   result_col38[30] <= result_col38[29];
   result_col38[31] <= result_col38[30];
   result_col38[32] <= result_col38[31];
   result_col38[33] <= result_col38[32];
   result_col38[34] <= result_col38[33];
   result_col38[35] <= result_col38[34];
   result_col38[36] <= result_col38[35];
   result_col38[37] <= result_col38[36];
   result_col38[38] <= result_col38[37];
   result_col38[39] <= result_col38[38];
   result_col38[40] <= result_col38[39];
   result_col38[41] <= result_col38[40];
   result_col38[42] <= result_col38[41];
   result_col38[43] <= result_col38[42];
   result_col38[44] <= result_col38[43];
   result_col38[45] <= result_col38[44];
   result_col38[46] <= result_col38[45];
   result_col38[47] <= result_col38[46];
   result_col38[48] <= result_col38[47];
   result_col38[49] <= result_col38[48];
   result_col38[50] <= result_col38[49];
   result_col38[51] <= result_col38[50];
   result_col38[52] <= result_col38[51];
   result_col38[53] <= result_col38[52];
   result_col38[54] <= result_col38[53];
   result_col38[55] <= result_col38[54];
   result_col38[56] <= result_col38[55];
   result_col38[57] <= result_col38[56];
   result_col38[58] <= result_col38[57];
   result_col38[59] <= result_col38[58];
   result_col38[60] <= result_col38[59];
   result_col38[61] <= result_col38[60];
   result_col38[62] <= result_col38[61];
   result_col38[63] <= result_col38[62];
   result_col38[64] <= result_col38[63];
   result_col38[65] <= result_col38[64];
   result_col38[66] <= result_col38[65];
   result_col38[67] <= result_col38[66];
   result_col38[68] <= result_col38[67];
   result_col38[69] <= result_col38[68];
   result_col38[70] <= result_col38[69];
   result_col38[71] <= result_col38[70];
   result_col38[72] <= result_col38[71];
   result_col38[73] <= result_col38[72];
   result_col38[74] <= result_col38[73];
   result_col38[75] <= result_col38[74];
   result_col38[76] <= result_col38[75];
   result_col38[77] <= result_col38[76];
   result_col38[78] <= result_col38[77];
   result_col38[79] <= result_col38[78];
   result_col38[80] <= result_col38[79];
   result_col38[81] <= result_col38[80];
   result_col38[82] <= result_col38[81];
   result_col38[83] <= result_col38[82];
   result_col38[84] <= result_col38[83];
   result_col38[85] <= result_col38[84];
   result_col38[86] <= result_col38[85];
   result_col38[87] <= result_col38[86];
   result_col38[88] <= result_col38[87];
   result_col38[89] <= result_col38[88];
   result_col38[90] <= result_col38[89];
   result_col38[91] <= result_col38[90];
   result_col38[92] <= result_col38[91];
   result_col38[93] <= result_col38[92];
   result_col38[94] <= result_col38[93];
   result_col38[95] <= result_col38[94];
   result_col38[96] <= result_col38[95];
   result_col38[97] <= result_col38[96];
   result_col38[98] <= result_col38[97];
   result_col38[99] <= result_col38[98];
   result_col38[100] <= result_col38[99];
   result_col38[101] <= result_col38[100];
   result_col38[102] <= result_col38[101];
   result_col38[103] <= result_col38[102];
   result_col38[104] <= result_col38[103];
   result_col38[105] <= result_col38[104];
   result_col38[106] <= result_col38[105];
   result_col38[107] <= result_col38[106];
   result_col38[108] <= result_col38[107];
   result_col38[109] <= result_col38[108];
   result_col38[110] <= result_col38[109];
   result_col38[111] <= result_col38[110];
   result_col38[112] <= result_col38[111];
   result_col38[113] <= result_col38[112];
   result_col38[114] <= result_col38[113];
   result_col38[115] <= result_col38[114];
   result_col38[116] <= result_col38[115];
   result_col38[117] <= result_col38[116];
   result_col38[118] <= result_col38[117];
   result_col38[119] <= result_col38[118];
   result_col38[120] <= result_col38[119];
   result_col38[121] <= result_col38[120];
   result_col38[122] <= result_col38[121];
   result_col38[123] <= result_col38[122];
   result_col38[124] <= result_col38[123];
   result_col38[125] <= result_col38[124];
   result_col38[126] <= result_col38[125];
   result_col38[127] <= result_col38[126];
   result_col38[128] <= result_col38[127];

   result_col39[1] <= data_out_4_39;
   result_col39[2] <= result_col39[1];
   result_col39[3] <= result_col39[2];
   result_col39[4] <= result_col39[3];
   result_col39[5] <= result_col39[4];
   result_col39[6] <= result_col39[5];
   result_col39[7] <= result_col39[6];
   result_col39[8] <= result_col39[7];
   result_col39[9] <= result_col39[8];
   result_col39[10] <= result_col39[9];
   result_col39[11] <= result_col39[10];
   result_col39[12] <= result_col39[11];
   result_col39[13] <= result_col39[12];
   result_col39[14] <= result_col39[13];
   result_col39[15] <= result_col39[14];
   result_col39[16] <= result_col39[15];
   result_col39[17] <= result_col39[16];
   result_col39[18] <= result_col39[17];
   result_col39[19] <= result_col39[18];
   result_col39[20] <= result_col39[19];
   result_col39[21] <= result_col39[20];
   result_col39[22] <= result_col39[21];
   result_col39[23] <= result_col39[22];
   result_col39[24] <= result_col39[23];
   result_col39[25] <= result_col39[24];
   result_col39[26] <= result_col39[25];
   result_col39[27] <= result_col39[26];
   result_col39[28] <= result_col39[27];
   result_col39[29] <= result_col39[28];
   result_col39[30] <= result_col39[29];
   result_col39[31] <= result_col39[30];
   result_col39[32] <= result_col39[31];
   result_col39[33] <= result_col39[32];
   result_col39[34] <= result_col39[33];
   result_col39[35] <= result_col39[34];
   result_col39[36] <= result_col39[35];
   result_col39[37] <= result_col39[36];
   result_col39[38] <= result_col39[37];
   result_col39[39] <= result_col39[38];
   result_col39[40] <= result_col39[39];
   result_col39[41] <= result_col39[40];
   result_col39[42] <= result_col39[41];
   result_col39[43] <= result_col39[42];
   result_col39[44] <= result_col39[43];
   result_col39[45] <= result_col39[44];
   result_col39[46] <= result_col39[45];
   result_col39[47] <= result_col39[46];
   result_col39[48] <= result_col39[47];
   result_col39[49] <= result_col39[48];
   result_col39[50] <= result_col39[49];
   result_col39[51] <= result_col39[50];
   result_col39[52] <= result_col39[51];
   result_col39[53] <= result_col39[52];
   result_col39[54] <= result_col39[53];
   result_col39[55] <= result_col39[54];
   result_col39[56] <= result_col39[55];
   result_col39[57] <= result_col39[56];
   result_col39[58] <= result_col39[57];
   result_col39[59] <= result_col39[58];
   result_col39[60] <= result_col39[59];
   result_col39[61] <= result_col39[60];
   result_col39[62] <= result_col39[61];
   result_col39[63] <= result_col39[62];
   result_col39[64] <= result_col39[63];
   result_col39[65] <= result_col39[64];
   result_col39[66] <= result_col39[65];
   result_col39[67] <= result_col39[66];
   result_col39[68] <= result_col39[67];
   result_col39[69] <= result_col39[68];
   result_col39[70] <= result_col39[69];
   result_col39[71] <= result_col39[70];
   result_col39[72] <= result_col39[71];
   result_col39[73] <= result_col39[72];
   result_col39[74] <= result_col39[73];
   result_col39[75] <= result_col39[74];
   result_col39[76] <= result_col39[75];
   result_col39[77] <= result_col39[76];
   result_col39[78] <= result_col39[77];
   result_col39[79] <= result_col39[78];
   result_col39[80] <= result_col39[79];
   result_col39[81] <= result_col39[80];
   result_col39[82] <= result_col39[81];
   result_col39[83] <= result_col39[82];
   result_col39[84] <= result_col39[83];
   result_col39[85] <= result_col39[84];
   result_col39[86] <= result_col39[85];
   result_col39[87] <= result_col39[86];
   result_col39[88] <= result_col39[87];
   result_col39[89] <= result_col39[88];
   result_col39[90] <= result_col39[89];
   result_col39[91] <= result_col39[90];
   result_col39[92] <= result_col39[91];
   result_col39[93] <= result_col39[92];
   result_col39[94] <= result_col39[93];
   result_col39[95] <= result_col39[94];
   result_col39[96] <= result_col39[95];
   result_col39[97] <= result_col39[96];
   result_col39[98] <= result_col39[97];
   result_col39[99] <= result_col39[98];
   result_col39[100] <= result_col39[99];
   result_col39[101] <= result_col39[100];
   result_col39[102] <= result_col39[101];
   result_col39[103] <= result_col39[102];
   result_col39[104] <= result_col39[103];
   result_col39[105] <= result_col39[104];
   result_col39[106] <= result_col39[105];
   result_col39[107] <= result_col39[106];
   result_col39[108] <= result_col39[107];
   result_col39[109] <= result_col39[108];
   result_col39[110] <= result_col39[109];
   result_col39[111] <= result_col39[110];
   result_col39[112] <= result_col39[111];
   result_col39[113] <= result_col39[112];
   result_col39[114] <= result_col39[113];
   result_col39[115] <= result_col39[114];
   result_col39[116] <= result_col39[115];
   result_col39[117] <= result_col39[116];
   result_col39[118] <= result_col39[117];
   result_col39[119] <= result_col39[118];
   result_col39[120] <= result_col39[119];
   result_col39[121] <= result_col39[120];
   result_col39[122] <= result_col39[121];
   result_col39[123] <= result_col39[122];
   result_col39[124] <= result_col39[123];
   result_col39[125] <= result_col39[124];
   result_col39[126] <= result_col39[125];
   result_col39[127] <= result_col39[126];

   result_col40[1] <= data_out_4_40;
   result_col40[2] <= result_col40[1];
   result_col40[3] <= result_col40[2];
   result_col40[4] <= result_col40[3];
   result_col40[5] <= result_col40[4];
   result_col40[6] <= result_col40[5];
   result_col40[7] <= result_col40[6];
   result_col40[8] <= result_col40[7];
   result_col40[9] <= result_col40[8];
   result_col40[10] <= result_col40[9];
   result_col40[11] <= result_col40[10];
   result_col40[12] <= result_col40[11];
   result_col40[13] <= result_col40[12];
   result_col40[14] <= result_col40[13];
   result_col40[15] <= result_col40[14];
   result_col40[16] <= result_col40[15];
   result_col40[17] <= result_col40[16];
   result_col40[18] <= result_col40[17];
   result_col40[19] <= result_col40[18];
   result_col40[20] <= result_col40[19];
   result_col40[21] <= result_col40[20];
   result_col40[22] <= result_col40[21];
   result_col40[23] <= result_col40[22];
   result_col40[24] <= result_col40[23];
   result_col40[25] <= result_col40[24];
   result_col40[26] <= result_col40[25];
   result_col40[27] <= result_col40[26];
   result_col40[28] <= result_col40[27];
   result_col40[29] <= result_col40[28];
   result_col40[30] <= result_col40[29];
   result_col40[31] <= result_col40[30];
   result_col40[32] <= result_col40[31];
   result_col40[33] <= result_col40[32];
   result_col40[34] <= result_col40[33];
   result_col40[35] <= result_col40[34];
   result_col40[36] <= result_col40[35];
   result_col40[37] <= result_col40[36];
   result_col40[38] <= result_col40[37];
   result_col40[39] <= result_col40[38];
   result_col40[40] <= result_col40[39];
   result_col40[41] <= result_col40[40];
   result_col40[42] <= result_col40[41];
   result_col40[43] <= result_col40[42];
   result_col40[44] <= result_col40[43];
   result_col40[45] <= result_col40[44];
   result_col40[46] <= result_col40[45];
   result_col40[47] <= result_col40[46];
   result_col40[48] <= result_col40[47];
   result_col40[49] <= result_col40[48];
   result_col40[50] <= result_col40[49];
   result_col40[51] <= result_col40[50];
   result_col40[52] <= result_col40[51];
   result_col40[53] <= result_col40[52];
   result_col40[54] <= result_col40[53];
   result_col40[55] <= result_col40[54];
   result_col40[56] <= result_col40[55];
   result_col40[57] <= result_col40[56];
   result_col40[58] <= result_col40[57];
   result_col40[59] <= result_col40[58];
   result_col40[60] <= result_col40[59];
   result_col40[61] <= result_col40[60];
   result_col40[62] <= result_col40[61];
   result_col40[63] <= result_col40[62];
   result_col40[64] <= result_col40[63];
   result_col40[65] <= result_col40[64];
   result_col40[66] <= result_col40[65];
   result_col40[67] <= result_col40[66];
   result_col40[68] <= result_col40[67];
   result_col40[69] <= result_col40[68];
   result_col40[70] <= result_col40[69];
   result_col40[71] <= result_col40[70];
   result_col40[72] <= result_col40[71];
   result_col40[73] <= result_col40[72];
   result_col40[74] <= result_col40[73];
   result_col40[75] <= result_col40[74];
   result_col40[76] <= result_col40[75];
   result_col40[77] <= result_col40[76];
   result_col40[78] <= result_col40[77];
   result_col40[79] <= result_col40[78];
   result_col40[80] <= result_col40[79];
   result_col40[81] <= result_col40[80];
   result_col40[82] <= result_col40[81];
   result_col40[83] <= result_col40[82];
   result_col40[84] <= result_col40[83];
   result_col40[85] <= result_col40[84];
   result_col40[86] <= result_col40[85];
   result_col40[87] <= result_col40[86];
   result_col40[88] <= result_col40[87];
   result_col40[89] <= result_col40[88];
   result_col40[90] <= result_col40[89];
   result_col40[91] <= result_col40[90];
   result_col40[92] <= result_col40[91];
   result_col40[93] <= result_col40[92];
   result_col40[94] <= result_col40[93];
   result_col40[95] <= result_col40[94];
   result_col40[96] <= result_col40[95];
   result_col40[97] <= result_col40[96];
   result_col40[98] <= result_col40[97];
   result_col40[99] <= result_col40[98];
   result_col40[100] <= result_col40[99];
   result_col40[101] <= result_col40[100];
   result_col40[102] <= result_col40[101];
   result_col40[103] <= result_col40[102];
   result_col40[104] <= result_col40[103];
   result_col40[105] <= result_col40[104];
   result_col40[106] <= result_col40[105];
   result_col40[107] <= result_col40[106];
   result_col40[108] <= result_col40[107];
   result_col40[109] <= result_col40[108];
   result_col40[110] <= result_col40[109];
   result_col40[111] <= result_col40[110];
   result_col40[112] <= result_col40[111];
   result_col40[113] <= result_col40[112];
   result_col40[114] <= result_col40[113];
   result_col40[115] <= result_col40[114];
   result_col40[116] <= result_col40[115];
   result_col40[117] <= result_col40[116];
   result_col40[118] <= result_col40[117];
   result_col40[119] <= result_col40[118];
   result_col40[120] <= result_col40[119];
   result_col40[121] <= result_col40[120];
   result_col40[122] <= result_col40[121];
   result_col40[123] <= result_col40[122];
   result_col40[124] <= result_col40[123];
   result_col40[125] <= result_col40[124];
   result_col40[126] <= result_col40[125];

   result_col41[1] <= data_out_4_41;
   result_col41[2] <= result_col41[1];
   result_col41[3] <= result_col41[2];
   result_col41[4] <= result_col41[3];
   result_col41[5] <= result_col41[4];
   result_col41[6] <= result_col41[5];
   result_col41[7] <= result_col41[6];
   result_col41[8] <= result_col41[7];
   result_col41[9] <= result_col41[8];
   result_col41[10] <= result_col41[9];
   result_col41[11] <= result_col41[10];
   result_col41[12] <= result_col41[11];
   result_col41[13] <= result_col41[12];
   result_col41[14] <= result_col41[13];
   result_col41[15] <= result_col41[14];
   result_col41[16] <= result_col41[15];
   result_col41[17] <= result_col41[16];
   result_col41[18] <= result_col41[17];
   result_col41[19] <= result_col41[18];
   result_col41[20] <= result_col41[19];
   result_col41[21] <= result_col41[20];
   result_col41[22] <= result_col41[21];
   result_col41[23] <= result_col41[22];
   result_col41[24] <= result_col41[23];
   result_col41[25] <= result_col41[24];
   result_col41[26] <= result_col41[25];
   result_col41[27] <= result_col41[26];
   result_col41[28] <= result_col41[27];
   result_col41[29] <= result_col41[28];
   result_col41[30] <= result_col41[29];
   result_col41[31] <= result_col41[30];
   result_col41[32] <= result_col41[31];
   result_col41[33] <= result_col41[32];
   result_col41[34] <= result_col41[33];
   result_col41[35] <= result_col41[34];
   result_col41[36] <= result_col41[35];
   result_col41[37] <= result_col41[36];
   result_col41[38] <= result_col41[37];
   result_col41[39] <= result_col41[38];
   result_col41[40] <= result_col41[39];
   result_col41[41] <= result_col41[40];
   result_col41[42] <= result_col41[41];
   result_col41[43] <= result_col41[42];
   result_col41[44] <= result_col41[43];
   result_col41[45] <= result_col41[44];
   result_col41[46] <= result_col41[45];
   result_col41[47] <= result_col41[46];
   result_col41[48] <= result_col41[47];
   result_col41[49] <= result_col41[48];
   result_col41[50] <= result_col41[49];
   result_col41[51] <= result_col41[50];
   result_col41[52] <= result_col41[51];
   result_col41[53] <= result_col41[52];
   result_col41[54] <= result_col41[53];
   result_col41[55] <= result_col41[54];
   result_col41[56] <= result_col41[55];
   result_col41[57] <= result_col41[56];
   result_col41[58] <= result_col41[57];
   result_col41[59] <= result_col41[58];
   result_col41[60] <= result_col41[59];
   result_col41[61] <= result_col41[60];
   result_col41[62] <= result_col41[61];
   result_col41[63] <= result_col41[62];
   result_col41[64] <= result_col41[63];
   result_col41[65] <= result_col41[64];
   result_col41[66] <= result_col41[65];
   result_col41[67] <= result_col41[66];
   result_col41[68] <= result_col41[67];
   result_col41[69] <= result_col41[68];
   result_col41[70] <= result_col41[69];
   result_col41[71] <= result_col41[70];
   result_col41[72] <= result_col41[71];
   result_col41[73] <= result_col41[72];
   result_col41[74] <= result_col41[73];
   result_col41[75] <= result_col41[74];
   result_col41[76] <= result_col41[75];
   result_col41[77] <= result_col41[76];
   result_col41[78] <= result_col41[77];
   result_col41[79] <= result_col41[78];
   result_col41[80] <= result_col41[79];
   result_col41[81] <= result_col41[80];
   result_col41[82] <= result_col41[81];
   result_col41[83] <= result_col41[82];
   result_col41[84] <= result_col41[83];
   result_col41[85] <= result_col41[84];
   result_col41[86] <= result_col41[85];
   result_col41[87] <= result_col41[86];
   result_col41[88] <= result_col41[87];
   result_col41[89] <= result_col41[88];
   result_col41[90] <= result_col41[89];
   result_col41[91] <= result_col41[90];
   result_col41[92] <= result_col41[91];
   result_col41[93] <= result_col41[92];
   result_col41[94] <= result_col41[93];
   result_col41[95] <= result_col41[94];
   result_col41[96] <= result_col41[95];
   result_col41[97] <= result_col41[96];
   result_col41[98] <= result_col41[97];
   result_col41[99] <= result_col41[98];
   result_col41[100] <= result_col41[99];
   result_col41[101] <= result_col41[100];
   result_col41[102] <= result_col41[101];
   result_col41[103] <= result_col41[102];
   result_col41[104] <= result_col41[103];
   result_col41[105] <= result_col41[104];
   result_col41[106] <= result_col41[105];
   result_col41[107] <= result_col41[106];
   result_col41[108] <= result_col41[107];
   result_col41[109] <= result_col41[108];
   result_col41[110] <= result_col41[109];
   result_col41[111] <= result_col41[110];
   result_col41[112] <= result_col41[111];
   result_col41[113] <= result_col41[112];
   result_col41[114] <= result_col41[113];
   result_col41[115] <= result_col41[114];
   result_col41[116] <= result_col41[115];
   result_col41[117] <= result_col41[116];
   result_col41[118] <= result_col41[117];
   result_col41[119] <= result_col41[118];
   result_col41[120] <= result_col41[119];
   result_col41[121] <= result_col41[120];
   result_col41[122] <= result_col41[121];
   result_col41[123] <= result_col41[122];
   result_col41[124] <= result_col41[123];
   result_col41[125] <= result_col41[124];

   result_col42[1] <= data_out_4_42;
   result_col42[2] <= result_col42[1];
   result_col42[3] <= result_col42[2];
   result_col42[4] <= result_col42[3];
   result_col42[5] <= result_col42[4];
   result_col42[6] <= result_col42[5];
   result_col42[7] <= result_col42[6];
   result_col42[8] <= result_col42[7];
   result_col42[9] <= result_col42[8];
   result_col42[10] <= result_col42[9];
   result_col42[11] <= result_col42[10];
   result_col42[12] <= result_col42[11];
   result_col42[13] <= result_col42[12];
   result_col42[14] <= result_col42[13];
   result_col42[15] <= result_col42[14];
   result_col42[16] <= result_col42[15];
   result_col42[17] <= result_col42[16];
   result_col42[18] <= result_col42[17];
   result_col42[19] <= result_col42[18];
   result_col42[20] <= result_col42[19];
   result_col42[21] <= result_col42[20];
   result_col42[22] <= result_col42[21];
   result_col42[23] <= result_col42[22];
   result_col42[24] <= result_col42[23];
   result_col42[25] <= result_col42[24];
   result_col42[26] <= result_col42[25];
   result_col42[27] <= result_col42[26];
   result_col42[28] <= result_col42[27];
   result_col42[29] <= result_col42[28];
   result_col42[30] <= result_col42[29];
   result_col42[31] <= result_col42[30];
   result_col42[32] <= result_col42[31];
   result_col42[33] <= result_col42[32];
   result_col42[34] <= result_col42[33];
   result_col42[35] <= result_col42[34];
   result_col42[36] <= result_col42[35];
   result_col42[37] <= result_col42[36];
   result_col42[38] <= result_col42[37];
   result_col42[39] <= result_col42[38];
   result_col42[40] <= result_col42[39];
   result_col42[41] <= result_col42[40];
   result_col42[42] <= result_col42[41];
   result_col42[43] <= result_col42[42];
   result_col42[44] <= result_col42[43];
   result_col42[45] <= result_col42[44];
   result_col42[46] <= result_col42[45];
   result_col42[47] <= result_col42[46];
   result_col42[48] <= result_col42[47];
   result_col42[49] <= result_col42[48];
   result_col42[50] <= result_col42[49];
   result_col42[51] <= result_col42[50];
   result_col42[52] <= result_col42[51];
   result_col42[53] <= result_col42[52];
   result_col42[54] <= result_col42[53];
   result_col42[55] <= result_col42[54];
   result_col42[56] <= result_col42[55];
   result_col42[57] <= result_col42[56];
   result_col42[58] <= result_col42[57];
   result_col42[59] <= result_col42[58];
   result_col42[60] <= result_col42[59];
   result_col42[61] <= result_col42[60];
   result_col42[62] <= result_col42[61];
   result_col42[63] <= result_col42[62];
   result_col42[64] <= result_col42[63];
   result_col42[65] <= result_col42[64];
   result_col42[66] <= result_col42[65];
   result_col42[67] <= result_col42[66];
   result_col42[68] <= result_col42[67];
   result_col42[69] <= result_col42[68];
   result_col42[70] <= result_col42[69];
   result_col42[71] <= result_col42[70];
   result_col42[72] <= result_col42[71];
   result_col42[73] <= result_col42[72];
   result_col42[74] <= result_col42[73];
   result_col42[75] <= result_col42[74];
   result_col42[76] <= result_col42[75];
   result_col42[77] <= result_col42[76];
   result_col42[78] <= result_col42[77];
   result_col42[79] <= result_col42[78];
   result_col42[80] <= result_col42[79];
   result_col42[81] <= result_col42[80];
   result_col42[82] <= result_col42[81];
   result_col42[83] <= result_col42[82];
   result_col42[84] <= result_col42[83];
   result_col42[85] <= result_col42[84];
   result_col42[86] <= result_col42[85];
   result_col42[87] <= result_col42[86];
   result_col42[88] <= result_col42[87];
   result_col42[89] <= result_col42[88];
   result_col42[90] <= result_col42[89];
   result_col42[91] <= result_col42[90];
   result_col42[92] <= result_col42[91];
   result_col42[93] <= result_col42[92];
   result_col42[94] <= result_col42[93];
   result_col42[95] <= result_col42[94];
   result_col42[96] <= result_col42[95];
   result_col42[97] <= result_col42[96];
   result_col42[98] <= result_col42[97];
   result_col42[99] <= result_col42[98];
   result_col42[100] <= result_col42[99];
   result_col42[101] <= result_col42[100];
   result_col42[102] <= result_col42[101];
   result_col42[103] <= result_col42[102];
   result_col42[104] <= result_col42[103];
   result_col42[105] <= result_col42[104];
   result_col42[106] <= result_col42[105];
   result_col42[107] <= result_col42[106];
   result_col42[108] <= result_col42[107];
   result_col42[109] <= result_col42[108];
   result_col42[110] <= result_col42[109];
   result_col42[111] <= result_col42[110];
   result_col42[112] <= result_col42[111];
   result_col42[113] <= result_col42[112];
   result_col42[114] <= result_col42[113];
   result_col42[115] <= result_col42[114];
   result_col42[116] <= result_col42[115];
   result_col42[117] <= result_col42[116];
   result_col42[118] <= result_col42[117];
   result_col42[119] <= result_col42[118];
   result_col42[120] <= result_col42[119];
   result_col42[121] <= result_col42[120];
   result_col42[122] <= result_col42[121];
   result_col42[123] <= result_col42[122];
   result_col42[124] <= result_col42[123];

   result_col43[1] <= data_out_4_43;
   result_col43[2] <= result_col43[1];
   result_col43[3] <= result_col43[2];
   result_col43[4] <= result_col43[3];
   result_col43[5] <= result_col43[4];
   result_col43[6] <= result_col43[5];
   result_col43[7] <= result_col43[6];
   result_col43[8] <= result_col43[7];
   result_col43[9] <= result_col43[8];
   result_col43[10] <= result_col43[9];
   result_col43[11] <= result_col43[10];
   result_col43[12] <= result_col43[11];
   result_col43[13] <= result_col43[12];
   result_col43[14] <= result_col43[13];
   result_col43[15] <= result_col43[14];
   result_col43[16] <= result_col43[15];
   result_col43[17] <= result_col43[16];
   result_col43[18] <= result_col43[17];
   result_col43[19] <= result_col43[18];
   result_col43[20] <= result_col43[19];
   result_col43[21] <= result_col43[20];
   result_col43[22] <= result_col43[21];
   result_col43[23] <= result_col43[22];
   result_col43[24] <= result_col43[23];
   result_col43[25] <= result_col43[24];
   result_col43[26] <= result_col43[25];
   result_col43[27] <= result_col43[26];
   result_col43[28] <= result_col43[27];
   result_col43[29] <= result_col43[28];
   result_col43[30] <= result_col43[29];
   result_col43[31] <= result_col43[30];
   result_col43[32] <= result_col43[31];
   result_col43[33] <= result_col43[32];
   result_col43[34] <= result_col43[33];
   result_col43[35] <= result_col43[34];
   result_col43[36] <= result_col43[35];
   result_col43[37] <= result_col43[36];
   result_col43[38] <= result_col43[37];
   result_col43[39] <= result_col43[38];
   result_col43[40] <= result_col43[39];
   result_col43[41] <= result_col43[40];
   result_col43[42] <= result_col43[41];
   result_col43[43] <= result_col43[42];
   result_col43[44] <= result_col43[43];
   result_col43[45] <= result_col43[44];
   result_col43[46] <= result_col43[45];
   result_col43[47] <= result_col43[46];
   result_col43[48] <= result_col43[47];
   result_col43[49] <= result_col43[48];
   result_col43[50] <= result_col43[49];
   result_col43[51] <= result_col43[50];
   result_col43[52] <= result_col43[51];
   result_col43[53] <= result_col43[52];
   result_col43[54] <= result_col43[53];
   result_col43[55] <= result_col43[54];
   result_col43[56] <= result_col43[55];
   result_col43[57] <= result_col43[56];
   result_col43[58] <= result_col43[57];
   result_col43[59] <= result_col43[58];
   result_col43[60] <= result_col43[59];
   result_col43[61] <= result_col43[60];
   result_col43[62] <= result_col43[61];
   result_col43[63] <= result_col43[62];
   result_col43[64] <= result_col43[63];
   result_col43[65] <= result_col43[64];
   result_col43[66] <= result_col43[65];
   result_col43[67] <= result_col43[66];
   result_col43[68] <= result_col43[67];
   result_col43[69] <= result_col43[68];
   result_col43[70] <= result_col43[69];
   result_col43[71] <= result_col43[70];
   result_col43[72] <= result_col43[71];
   result_col43[73] <= result_col43[72];
   result_col43[74] <= result_col43[73];
   result_col43[75] <= result_col43[74];
   result_col43[76] <= result_col43[75];
   result_col43[77] <= result_col43[76];
   result_col43[78] <= result_col43[77];
   result_col43[79] <= result_col43[78];
   result_col43[80] <= result_col43[79];
   result_col43[81] <= result_col43[80];
   result_col43[82] <= result_col43[81];
   result_col43[83] <= result_col43[82];
   result_col43[84] <= result_col43[83];
   result_col43[85] <= result_col43[84];
   result_col43[86] <= result_col43[85];
   result_col43[87] <= result_col43[86];
   result_col43[88] <= result_col43[87];
   result_col43[89] <= result_col43[88];
   result_col43[90] <= result_col43[89];
   result_col43[91] <= result_col43[90];
   result_col43[92] <= result_col43[91];
   result_col43[93] <= result_col43[92];
   result_col43[94] <= result_col43[93];
   result_col43[95] <= result_col43[94];
   result_col43[96] <= result_col43[95];
   result_col43[97] <= result_col43[96];
   result_col43[98] <= result_col43[97];
   result_col43[99] <= result_col43[98];
   result_col43[100] <= result_col43[99];
   result_col43[101] <= result_col43[100];
   result_col43[102] <= result_col43[101];
   result_col43[103] <= result_col43[102];
   result_col43[104] <= result_col43[103];
   result_col43[105] <= result_col43[104];
   result_col43[106] <= result_col43[105];
   result_col43[107] <= result_col43[106];
   result_col43[108] <= result_col43[107];
   result_col43[109] <= result_col43[108];
   result_col43[110] <= result_col43[109];
   result_col43[111] <= result_col43[110];
   result_col43[112] <= result_col43[111];
   result_col43[113] <= result_col43[112];
   result_col43[114] <= result_col43[113];
   result_col43[115] <= result_col43[114];
   result_col43[116] <= result_col43[115];
   result_col43[117] <= result_col43[116];
   result_col43[118] <= result_col43[117];
   result_col43[119] <= result_col43[118];
   result_col43[120] <= result_col43[119];
   result_col43[121] <= result_col43[120];
   result_col43[122] <= result_col43[121];
   result_col43[123] <= result_col43[122];

   result_col44[1] <= data_out_4_44;
   result_col44[2] <= result_col44[1];
   result_col44[3] <= result_col44[2];
   result_col44[4] <= result_col44[3];
   result_col44[5] <= result_col44[4];
   result_col44[6] <= result_col44[5];
   result_col44[7] <= result_col44[6];
   result_col44[8] <= result_col44[7];
   result_col44[9] <= result_col44[8];
   result_col44[10] <= result_col44[9];
   result_col44[11] <= result_col44[10];
   result_col44[12] <= result_col44[11];
   result_col44[13] <= result_col44[12];
   result_col44[14] <= result_col44[13];
   result_col44[15] <= result_col44[14];
   result_col44[16] <= result_col44[15];
   result_col44[17] <= result_col44[16];
   result_col44[18] <= result_col44[17];
   result_col44[19] <= result_col44[18];
   result_col44[20] <= result_col44[19];
   result_col44[21] <= result_col44[20];
   result_col44[22] <= result_col44[21];
   result_col44[23] <= result_col44[22];
   result_col44[24] <= result_col44[23];
   result_col44[25] <= result_col44[24];
   result_col44[26] <= result_col44[25];
   result_col44[27] <= result_col44[26];
   result_col44[28] <= result_col44[27];
   result_col44[29] <= result_col44[28];
   result_col44[30] <= result_col44[29];
   result_col44[31] <= result_col44[30];
   result_col44[32] <= result_col44[31];
   result_col44[33] <= result_col44[32];
   result_col44[34] <= result_col44[33];
   result_col44[35] <= result_col44[34];
   result_col44[36] <= result_col44[35];
   result_col44[37] <= result_col44[36];
   result_col44[38] <= result_col44[37];
   result_col44[39] <= result_col44[38];
   result_col44[40] <= result_col44[39];
   result_col44[41] <= result_col44[40];
   result_col44[42] <= result_col44[41];
   result_col44[43] <= result_col44[42];
   result_col44[44] <= result_col44[43];
   result_col44[45] <= result_col44[44];
   result_col44[46] <= result_col44[45];
   result_col44[47] <= result_col44[46];
   result_col44[48] <= result_col44[47];
   result_col44[49] <= result_col44[48];
   result_col44[50] <= result_col44[49];
   result_col44[51] <= result_col44[50];
   result_col44[52] <= result_col44[51];
   result_col44[53] <= result_col44[52];
   result_col44[54] <= result_col44[53];
   result_col44[55] <= result_col44[54];
   result_col44[56] <= result_col44[55];
   result_col44[57] <= result_col44[56];
   result_col44[58] <= result_col44[57];
   result_col44[59] <= result_col44[58];
   result_col44[60] <= result_col44[59];
   result_col44[61] <= result_col44[60];
   result_col44[62] <= result_col44[61];
   result_col44[63] <= result_col44[62];
   result_col44[64] <= result_col44[63];
   result_col44[65] <= result_col44[64];
   result_col44[66] <= result_col44[65];
   result_col44[67] <= result_col44[66];
   result_col44[68] <= result_col44[67];
   result_col44[69] <= result_col44[68];
   result_col44[70] <= result_col44[69];
   result_col44[71] <= result_col44[70];
   result_col44[72] <= result_col44[71];
   result_col44[73] <= result_col44[72];
   result_col44[74] <= result_col44[73];
   result_col44[75] <= result_col44[74];
   result_col44[76] <= result_col44[75];
   result_col44[77] <= result_col44[76];
   result_col44[78] <= result_col44[77];
   result_col44[79] <= result_col44[78];
   result_col44[80] <= result_col44[79];
   result_col44[81] <= result_col44[80];
   result_col44[82] <= result_col44[81];
   result_col44[83] <= result_col44[82];
   result_col44[84] <= result_col44[83];
   result_col44[85] <= result_col44[84];
   result_col44[86] <= result_col44[85];
   result_col44[87] <= result_col44[86];
   result_col44[88] <= result_col44[87];
   result_col44[89] <= result_col44[88];
   result_col44[90] <= result_col44[89];
   result_col44[91] <= result_col44[90];
   result_col44[92] <= result_col44[91];
   result_col44[93] <= result_col44[92];
   result_col44[94] <= result_col44[93];
   result_col44[95] <= result_col44[94];
   result_col44[96] <= result_col44[95];
   result_col44[97] <= result_col44[96];
   result_col44[98] <= result_col44[97];
   result_col44[99] <= result_col44[98];
   result_col44[100] <= result_col44[99];
   result_col44[101] <= result_col44[100];
   result_col44[102] <= result_col44[101];
   result_col44[103] <= result_col44[102];
   result_col44[104] <= result_col44[103];
   result_col44[105] <= result_col44[104];
   result_col44[106] <= result_col44[105];
   result_col44[107] <= result_col44[106];
   result_col44[108] <= result_col44[107];
   result_col44[109] <= result_col44[108];
   result_col44[110] <= result_col44[109];
   result_col44[111] <= result_col44[110];
   result_col44[112] <= result_col44[111];
   result_col44[113] <= result_col44[112];
   result_col44[114] <= result_col44[113];
   result_col44[115] <= result_col44[114];
   result_col44[116] <= result_col44[115];
   result_col44[117] <= result_col44[116];
   result_col44[118] <= result_col44[117];
   result_col44[119] <= result_col44[118];
   result_col44[120] <= result_col44[119];
   result_col44[121] <= result_col44[120];
   result_col44[122] <= result_col44[121];

   result_col45[1] <= data_out_4_45;
   result_col45[2] <= result_col45[1];
   result_col45[3] <= result_col45[2];
   result_col45[4] <= result_col45[3];
   result_col45[5] <= result_col45[4];
   result_col45[6] <= result_col45[5];
   result_col45[7] <= result_col45[6];
   result_col45[8] <= result_col45[7];
   result_col45[9] <= result_col45[8];
   result_col45[10] <= result_col45[9];
   result_col45[11] <= result_col45[10];
   result_col45[12] <= result_col45[11];
   result_col45[13] <= result_col45[12];
   result_col45[14] <= result_col45[13];
   result_col45[15] <= result_col45[14];
   result_col45[16] <= result_col45[15];
   result_col45[17] <= result_col45[16];
   result_col45[18] <= result_col45[17];
   result_col45[19] <= result_col45[18];
   result_col45[20] <= result_col45[19];
   result_col45[21] <= result_col45[20];
   result_col45[22] <= result_col45[21];
   result_col45[23] <= result_col45[22];
   result_col45[24] <= result_col45[23];
   result_col45[25] <= result_col45[24];
   result_col45[26] <= result_col45[25];
   result_col45[27] <= result_col45[26];
   result_col45[28] <= result_col45[27];
   result_col45[29] <= result_col45[28];
   result_col45[30] <= result_col45[29];
   result_col45[31] <= result_col45[30];
   result_col45[32] <= result_col45[31];
   result_col45[33] <= result_col45[32];
   result_col45[34] <= result_col45[33];
   result_col45[35] <= result_col45[34];
   result_col45[36] <= result_col45[35];
   result_col45[37] <= result_col45[36];
   result_col45[38] <= result_col45[37];
   result_col45[39] <= result_col45[38];
   result_col45[40] <= result_col45[39];
   result_col45[41] <= result_col45[40];
   result_col45[42] <= result_col45[41];
   result_col45[43] <= result_col45[42];
   result_col45[44] <= result_col45[43];
   result_col45[45] <= result_col45[44];
   result_col45[46] <= result_col45[45];
   result_col45[47] <= result_col45[46];
   result_col45[48] <= result_col45[47];
   result_col45[49] <= result_col45[48];
   result_col45[50] <= result_col45[49];
   result_col45[51] <= result_col45[50];
   result_col45[52] <= result_col45[51];
   result_col45[53] <= result_col45[52];
   result_col45[54] <= result_col45[53];
   result_col45[55] <= result_col45[54];
   result_col45[56] <= result_col45[55];
   result_col45[57] <= result_col45[56];
   result_col45[58] <= result_col45[57];
   result_col45[59] <= result_col45[58];
   result_col45[60] <= result_col45[59];
   result_col45[61] <= result_col45[60];
   result_col45[62] <= result_col45[61];
   result_col45[63] <= result_col45[62];
   result_col45[64] <= result_col45[63];
   result_col45[65] <= result_col45[64];
   result_col45[66] <= result_col45[65];
   result_col45[67] <= result_col45[66];
   result_col45[68] <= result_col45[67];
   result_col45[69] <= result_col45[68];
   result_col45[70] <= result_col45[69];
   result_col45[71] <= result_col45[70];
   result_col45[72] <= result_col45[71];
   result_col45[73] <= result_col45[72];
   result_col45[74] <= result_col45[73];
   result_col45[75] <= result_col45[74];
   result_col45[76] <= result_col45[75];
   result_col45[77] <= result_col45[76];
   result_col45[78] <= result_col45[77];
   result_col45[79] <= result_col45[78];
   result_col45[80] <= result_col45[79];
   result_col45[81] <= result_col45[80];
   result_col45[82] <= result_col45[81];
   result_col45[83] <= result_col45[82];
   result_col45[84] <= result_col45[83];
   result_col45[85] <= result_col45[84];
   result_col45[86] <= result_col45[85];
   result_col45[87] <= result_col45[86];
   result_col45[88] <= result_col45[87];
   result_col45[89] <= result_col45[88];
   result_col45[90] <= result_col45[89];
   result_col45[91] <= result_col45[90];
   result_col45[92] <= result_col45[91];
   result_col45[93] <= result_col45[92];
   result_col45[94] <= result_col45[93];
   result_col45[95] <= result_col45[94];
   result_col45[96] <= result_col45[95];
   result_col45[97] <= result_col45[96];
   result_col45[98] <= result_col45[97];
   result_col45[99] <= result_col45[98];
   result_col45[100] <= result_col45[99];
   result_col45[101] <= result_col45[100];
   result_col45[102] <= result_col45[101];
   result_col45[103] <= result_col45[102];
   result_col45[104] <= result_col45[103];
   result_col45[105] <= result_col45[104];
   result_col45[106] <= result_col45[105];
   result_col45[107] <= result_col45[106];
   result_col45[108] <= result_col45[107];
   result_col45[109] <= result_col45[108];
   result_col45[110] <= result_col45[109];
   result_col45[111] <= result_col45[110];
   result_col45[112] <= result_col45[111];
   result_col45[113] <= result_col45[112];
   result_col45[114] <= result_col45[113];
   result_col45[115] <= result_col45[114];
   result_col45[116] <= result_col45[115];
   result_col45[117] <= result_col45[116];
   result_col45[118] <= result_col45[117];
   result_col45[119] <= result_col45[118];
   result_col45[120] <= result_col45[119];
   result_col45[121] <= result_col45[120];

   result_col46[1] <= data_out_4_46;
   result_col46[2] <= result_col46[1];
   result_col46[3] <= result_col46[2];
   result_col46[4] <= result_col46[3];
   result_col46[5] <= result_col46[4];
   result_col46[6] <= result_col46[5];
   result_col46[7] <= result_col46[6];
   result_col46[8] <= result_col46[7];
   result_col46[9] <= result_col46[8];
   result_col46[10] <= result_col46[9];
   result_col46[11] <= result_col46[10];
   result_col46[12] <= result_col46[11];
   result_col46[13] <= result_col46[12];
   result_col46[14] <= result_col46[13];
   result_col46[15] <= result_col46[14];
   result_col46[16] <= result_col46[15];
   result_col46[17] <= result_col46[16];
   result_col46[18] <= result_col46[17];
   result_col46[19] <= result_col46[18];
   result_col46[20] <= result_col46[19];
   result_col46[21] <= result_col46[20];
   result_col46[22] <= result_col46[21];
   result_col46[23] <= result_col46[22];
   result_col46[24] <= result_col46[23];
   result_col46[25] <= result_col46[24];
   result_col46[26] <= result_col46[25];
   result_col46[27] <= result_col46[26];
   result_col46[28] <= result_col46[27];
   result_col46[29] <= result_col46[28];
   result_col46[30] <= result_col46[29];
   result_col46[31] <= result_col46[30];
   result_col46[32] <= result_col46[31];
   result_col46[33] <= result_col46[32];
   result_col46[34] <= result_col46[33];
   result_col46[35] <= result_col46[34];
   result_col46[36] <= result_col46[35];
   result_col46[37] <= result_col46[36];
   result_col46[38] <= result_col46[37];
   result_col46[39] <= result_col46[38];
   result_col46[40] <= result_col46[39];
   result_col46[41] <= result_col46[40];
   result_col46[42] <= result_col46[41];
   result_col46[43] <= result_col46[42];
   result_col46[44] <= result_col46[43];
   result_col46[45] <= result_col46[44];
   result_col46[46] <= result_col46[45];
   result_col46[47] <= result_col46[46];
   result_col46[48] <= result_col46[47];
   result_col46[49] <= result_col46[48];
   result_col46[50] <= result_col46[49];
   result_col46[51] <= result_col46[50];
   result_col46[52] <= result_col46[51];
   result_col46[53] <= result_col46[52];
   result_col46[54] <= result_col46[53];
   result_col46[55] <= result_col46[54];
   result_col46[56] <= result_col46[55];
   result_col46[57] <= result_col46[56];
   result_col46[58] <= result_col46[57];
   result_col46[59] <= result_col46[58];
   result_col46[60] <= result_col46[59];
   result_col46[61] <= result_col46[60];
   result_col46[62] <= result_col46[61];
   result_col46[63] <= result_col46[62];
   result_col46[64] <= result_col46[63];
   result_col46[65] <= result_col46[64];
   result_col46[66] <= result_col46[65];
   result_col46[67] <= result_col46[66];
   result_col46[68] <= result_col46[67];
   result_col46[69] <= result_col46[68];
   result_col46[70] <= result_col46[69];
   result_col46[71] <= result_col46[70];
   result_col46[72] <= result_col46[71];
   result_col46[73] <= result_col46[72];
   result_col46[74] <= result_col46[73];
   result_col46[75] <= result_col46[74];
   result_col46[76] <= result_col46[75];
   result_col46[77] <= result_col46[76];
   result_col46[78] <= result_col46[77];
   result_col46[79] <= result_col46[78];
   result_col46[80] <= result_col46[79];
   result_col46[81] <= result_col46[80];
   result_col46[82] <= result_col46[81];
   result_col46[83] <= result_col46[82];
   result_col46[84] <= result_col46[83];
   result_col46[85] <= result_col46[84];
   result_col46[86] <= result_col46[85];
   result_col46[87] <= result_col46[86];
   result_col46[88] <= result_col46[87];
   result_col46[89] <= result_col46[88];
   result_col46[90] <= result_col46[89];
   result_col46[91] <= result_col46[90];
   result_col46[92] <= result_col46[91];
   result_col46[93] <= result_col46[92];
   result_col46[94] <= result_col46[93];
   result_col46[95] <= result_col46[94];
   result_col46[96] <= result_col46[95];
   result_col46[97] <= result_col46[96];
   result_col46[98] <= result_col46[97];
   result_col46[99] <= result_col46[98];
   result_col46[100] <= result_col46[99];
   result_col46[101] <= result_col46[100];
   result_col46[102] <= result_col46[101];
   result_col46[103] <= result_col46[102];
   result_col46[104] <= result_col46[103];
   result_col46[105] <= result_col46[104];
   result_col46[106] <= result_col46[105];
   result_col46[107] <= result_col46[106];
   result_col46[108] <= result_col46[107];
   result_col46[109] <= result_col46[108];
   result_col46[110] <= result_col46[109];
   result_col46[111] <= result_col46[110];
   result_col46[112] <= result_col46[111];
   result_col46[113] <= result_col46[112];
   result_col46[114] <= result_col46[113];
   result_col46[115] <= result_col46[114];
   result_col46[116] <= result_col46[115];
   result_col46[117] <= result_col46[116];
   result_col46[118] <= result_col46[117];
   result_col46[119] <= result_col46[118];
   result_col46[120] <= result_col46[119];

   result_col47[1] <= data_out_4_47;
   result_col47[2] <= result_col47[1];
   result_col47[3] <= result_col47[2];
   result_col47[4] <= result_col47[3];
   result_col47[5] <= result_col47[4];
   result_col47[6] <= result_col47[5];
   result_col47[7] <= result_col47[6];
   result_col47[8] <= result_col47[7];
   result_col47[9] <= result_col47[8];
   result_col47[10] <= result_col47[9];
   result_col47[11] <= result_col47[10];
   result_col47[12] <= result_col47[11];
   result_col47[13] <= result_col47[12];
   result_col47[14] <= result_col47[13];
   result_col47[15] <= result_col47[14];
   result_col47[16] <= result_col47[15];
   result_col47[17] <= result_col47[16];
   result_col47[18] <= result_col47[17];
   result_col47[19] <= result_col47[18];
   result_col47[20] <= result_col47[19];
   result_col47[21] <= result_col47[20];
   result_col47[22] <= result_col47[21];
   result_col47[23] <= result_col47[22];
   result_col47[24] <= result_col47[23];
   result_col47[25] <= result_col47[24];
   result_col47[26] <= result_col47[25];
   result_col47[27] <= result_col47[26];
   result_col47[28] <= result_col47[27];
   result_col47[29] <= result_col47[28];
   result_col47[30] <= result_col47[29];
   result_col47[31] <= result_col47[30];
   result_col47[32] <= result_col47[31];
   result_col47[33] <= result_col47[32];
   result_col47[34] <= result_col47[33];
   result_col47[35] <= result_col47[34];
   result_col47[36] <= result_col47[35];
   result_col47[37] <= result_col47[36];
   result_col47[38] <= result_col47[37];
   result_col47[39] <= result_col47[38];
   result_col47[40] <= result_col47[39];
   result_col47[41] <= result_col47[40];
   result_col47[42] <= result_col47[41];
   result_col47[43] <= result_col47[42];
   result_col47[44] <= result_col47[43];
   result_col47[45] <= result_col47[44];
   result_col47[46] <= result_col47[45];
   result_col47[47] <= result_col47[46];
   result_col47[48] <= result_col47[47];
   result_col47[49] <= result_col47[48];
   result_col47[50] <= result_col47[49];
   result_col47[51] <= result_col47[50];
   result_col47[52] <= result_col47[51];
   result_col47[53] <= result_col47[52];
   result_col47[54] <= result_col47[53];
   result_col47[55] <= result_col47[54];
   result_col47[56] <= result_col47[55];
   result_col47[57] <= result_col47[56];
   result_col47[58] <= result_col47[57];
   result_col47[59] <= result_col47[58];
   result_col47[60] <= result_col47[59];
   result_col47[61] <= result_col47[60];
   result_col47[62] <= result_col47[61];
   result_col47[63] <= result_col47[62];
   result_col47[64] <= result_col47[63];
   result_col47[65] <= result_col47[64];
   result_col47[66] <= result_col47[65];
   result_col47[67] <= result_col47[66];
   result_col47[68] <= result_col47[67];
   result_col47[69] <= result_col47[68];
   result_col47[70] <= result_col47[69];
   result_col47[71] <= result_col47[70];
   result_col47[72] <= result_col47[71];
   result_col47[73] <= result_col47[72];
   result_col47[74] <= result_col47[73];
   result_col47[75] <= result_col47[74];
   result_col47[76] <= result_col47[75];
   result_col47[77] <= result_col47[76];
   result_col47[78] <= result_col47[77];
   result_col47[79] <= result_col47[78];
   result_col47[80] <= result_col47[79];
   result_col47[81] <= result_col47[80];
   result_col47[82] <= result_col47[81];
   result_col47[83] <= result_col47[82];
   result_col47[84] <= result_col47[83];
   result_col47[85] <= result_col47[84];
   result_col47[86] <= result_col47[85];
   result_col47[87] <= result_col47[86];
   result_col47[88] <= result_col47[87];
   result_col47[89] <= result_col47[88];
   result_col47[90] <= result_col47[89];
   result_col47[91] <= result_col47[90];
   result_col47[92] <= result_col47[91];
   result_col47[93] <= result_col47[92];
   result_col47[94] <= result_col47[93];
   result_col47[95] <= result_col47[94];
   result_col47[96] <= result_col47[95];
   result_col47[97] <= result_col47[96];
   result_col47[98] <= result_col47[97];
   result_col47[99] <= result_col47[98];
   result_col47[100] <= result_col47[99];
   result_col47[101] <= result_col47[100];
   result_col47[102] <= result_col47[101];
   result_col47[103] <= result_col47[102];
   result_col47[104] <= result_col47[103];
   result_col47[105] <= result_col47[104];
   result_col47[106] <= result_col47[105];
   result_col47[107] <= result_col47[106];
   result_col47[108] <= result_col47[107];
   result_col47[109] <= result_col47[108];
   result_col47[110] <= result_col47[109];
   result_col47[111] <= result_col47[110];
   result_col47[112] <= result_col47[111];
   result_col47[113] <= result_col47[112];
   result_col47[114] <= result_col47[113];
   result_col47[115] <= result_col47[114];
   result_col47[116] <= result_col47[115];
   result_col47[117] <= result_col47[116];
   result_col47[118] <= result_col47[117];
   result_col47[119] <= result_col47[118];

   result_col48[1] <= data_out_4_48;
   result_col48[2] <= result_col48[1];
   result_col48[3] <= result_col48[2];
   result_col48[4] <= result_col48[3];
   result_col48[5] <= result_col48[4];
   result_col48[6] <= result_col48[5];
   result_col48[7] <= result_col48[6];
   result_col48[8] <= result_col48[7];
   result_col48[9] <= result_col48[8];
   result_col48[10] <= result_col48[9];
   result_col48[11] <= result_col48[10];
   result_col48[12] <= result_col48[11];
   result_col48[13] <= result_col48[12];
   result_col48[14] <= result_col48[13];
   result_col48[15] <= result_col48[14];
   result_col48[16] <= result_col48[15];
   result_col48[17] <= result_col48[16];
   result_col48[18] <= result_col48[17];
   result_col48[19] <= result_col48[18];
   result_col48[20] <= result_col48[19];
   result_col48[21] <= result_col48[20];
   result_col48[22] <= result_col48[21];
   result_col48[23] <= result_col48[22];
   result_col48[24] <= result_col48[23];
   result_col48[25] <= result_col48[24];
   result_col48[26] <= result_col48[25];
   result_col48[27] <= result_col48[26];
   result_col48[28] <= result_col48[27];
   result_col48[29] <= result_col48[28];
   result_col48[30] <= result_col48[29];
   result_col48[31] <= result_col48[30];
   result_col48[32] <= result_col48[31];
   result_col48[33] <= result_col48[32];
   result_col48[34] <= result_col48[33];
   result_col48[35] <= result_col48[34];
   result_col48[36] <= result_col48[35];
   result_col48[37] <= result_col48[36];
   result_col48[38] <= result_col48[37];
   result_col48[39] <= result_col48[38];
   result_col48[40] <= result_col48[39];
   result_col48[41] <= result_col48[40];
   result_col48[42] <= result_col48[41];
   result_col48[43] <= result_col48[42];
   result_col48[44] <= result_col48[43];
   result_col48[45] <= result_col48[44];
   result_col48[46] <= result_col48[45];
   result_col48[47] <= result_col48[46];
   result_col48[48] <= result_col48[47];
   result_col48[49] <= result_col48[48];
   result_col48[50] <= result_col48[49];
   result_col48[51] <= result_col48[50];
   result_col48[52] <= result_col48[51];
   result_col48[53] <= result_col48[52];
   result_col48[54] <= result_col48[53];
   result_col48[55] <= result_col48[54];
   result_col48[56] <= result_col48[55];
   result_col48[57] <= result_col48[56];
   result_col48[58] <= result_col48[57];
   result_col48[59] <= result_col48[58];
   result_col48[60] <= result_col48[59];
   result_col48[61] <= result_col48[60];
   result_col48[62] <= result_col48[61];
   result_col48[63] <= result_col48[62];
   result_col48[64] <= result_col48[63];
   result_col48[65] <= result_col48[64];
   result_col48[66] <= result_col48[65];
   result_col48[67] <= result_col48[66];
   result_col48[68] <= result_col48[67];
   result_col48[69] <= result_col48[68];
   result_col48[70] <= result_col48[69];
   result_col48[71] <= result_col48[70];
   result_col48[72] <= result_col48[71];
   result_col48[73] <= result_col48[72];
   result_col48[74] <= result_col48[73];
   result_col48[75] <= result_col48[74];
   result_col48[76] <= result_col48[75];
   result_col48[77] <= result_col48[76];
   result_col48[78] <= result_col48[77];
   result_col48[79] <= result_col48[78];
   result_col48[80] <= result_col48[79];
   result_col48[81] <= result_col48[80];
   result_col48[82] <= result_col48[81];
   result_col48[83] <= result_col48[82];
   result_col48[84] <= result_col48[83];
   result_col48[85] <= result_col48[84];
   result_col48[86] <= result_col48[85];
   result_col48[87] <= result_col48[86];
   result_col48[88] <= result_col48[87];
   result_col48[89] <= result_col48[88];
   result_col48[90] <= result_col48[89];
   result_col48[91] <= result_col48[90];
   result_col48[92] <= result_col48[91];
   result_col48[93] <= result_col48[92];
   result_col48[94] <= result_col48[93];
   result_col48[95] <= result_col48[94];
   result_col48[96] <= result_col48[95];
   result_col48[97] <= result_col48[96];
   result_col48[98] <= result_col48[97];
   result_col48[99] <= result_col48[98];
   result_col48[100] <= result_col48[99];
   result_col48[101] <= result_col48[100];
   result_col48[102] <= result_col48[101];
   result_col48[103] <= result_col48[102];
   result_col48[104] <= result_col48[103];
   result_col48[105] <= result_col48[104];
   result_col48[106] <= result_col48[105];
   result_col48[107] <= result_col48[106];
   result_col48[108] <= result_col48[107];
   result_col48[109] <= result_col48[108];
   result_col48[110] <= result_col48[109];
   result_col48[111] <= result_col48[110];
   result_col48[112] <= result_col48[111];
   result_col48[113] <= result_col48[112];
   result_col48[114] <= result_col48[113];
   result_col48[115] <= result_col48[114];
   result_col48[116] <= result_col48[115];
   result_col48[117] <= result_col48[116];
   result_col48[118] <= result_col48[117];

   result_col49[1] <= data_out_4_49;
   result_col49[2] <= result_col49[1];
   result_col49[3] <= result_col49[2];
   result_col49[4] <= result_col49[3];
   result_col49[5] <= result_col49[4];
   result_col49[6] <= result_col49[5];
   result_col49[7] <= result_col49[6];
   result_col49[8] <= result_col49[7];
   result_col49[9] <= result_col49[8];
   result_col49[10] <= result_col49[9];
   result_col49[11] <= result_col49[10];
   result_col49[12] <= result_col49[11];
   result_col49[13] <= result_col49[12];
   result_col49[14] <= result_col49[13];
   result_col49[15] <= result_col49[14];
   result_col49[16] <= result_col49[15];
   result_col49[17] <= result_col49[16];
   result_col49[18] <= result_col49[17];
   result_col49[19] <= result_col49[18];
   result_col49[20] <= result_col49[19];
   result_col49[21] <= result_col49[20];
   result_col49[22] <= result_col49[21];
   result_col49[23] <= result_col49[22];
   result_col49[24] <= result_col49[23];
   result_col49[25] <= result_col49[24];
   result_col49[26] <= result_col49[25];
   result_col49[27] <= result_col49[26];
   result_col49[28] <= result_col49[27];
   result_col49[29] <= result_col49[28];
   result_col49[30] <= result_col49[29];
   result_col49[31] <= result_col49[30];
   result_col49[32] <= result_col49[31];
   result_col49[33] <= result_col49[32];
   result_col49[34] <= result_col49[33];
   result_col49[35] <= result_col49[34];
   result_col49[36] <= result_col49[35];
   result_col49[37] <= result_col49[36];
   result_col49[38] <= result_col49[37];
   result_col49[39] <= result_col49[38];
   result_col49[40] <= result_col49[39];
   result_col49[41] <= result_col49[40];
   result_col49[42] <= result_col49[41];
   result_col49[43] <= result_col49[42];
   result_col49[44] <= result_col49[43];
   result_col49[45] <= result_col49[44];
   result_col49[46] <= result_col49[45];
   result_col49[47] <= result_col49[46];
   result_col49[48] <= result_col49[47];
   result_col49[49] <= result_col49[48];
   result_col49[50] <= result_col49[49];
   result_col49[51] <= result_col49[50];
   result_col49[52] <= result_col49[51];
   result_col49[53] <= result_col49[52];
   result_col49[54] <= result_col49[53];
   result_col49[55] <= result_col49[54];
   result_col49[56] <= result_col49[55];
   result_col49[57] <= result_col49[56];
   result_col49[58] <= result_col49[57];
   result_col49[59] <= result_col49[58];
   result_col49[60] <= result_col49[59];
   result_col49[61] <= result_col49[60];
   result_col49[62] <= result_col49[61];
   result_col49[63] <= result_col49[62];
   result_col49[64] <= result_col49[63];
   result_col49[65] <= result_col49[64];
   result_col49[66] <= result_col49[65];
   result_col49[67] <= result_col49[66];
   result_col49[68] <= result_col49[67];
   result_col49[69] <= result_col49[68];
   result_col49[70] <= result_col49[69];
   result_col49[71] <= result_col49[70];
   result_col49[72] <= result_col49[71];
   result_col49[73] <= result_col49[72];
   result_col49[74] <= result_col49[73];
   result_col49[75] <= result_col49[74];
   result_col49[76] <= result_col49[75];
   result_col49[77] <= result_col49[76];
   result_col49[78] <= result_col49[77];
   result_col49[79] <= result_col49[78];
   result_col49[80] <= result_col49[79];
   result_col49[81] <= result_col49[80];
   result_col49[82] <= result_col49[81];
   result_col49[83] <= result_col49[82];
   result_col49[84] <= result_col49[83];
   result_col49[85] <= result_col49[84];
   result_col49[86] <= result_col49[85];
   result_col49[87] <= result_col49[86];
   result_col49[88] <= result_col49[87];
   result_col49[89] <= result_col49[88];
   result_col49[90] <= result_col49[89];
   result_col49[91] <= result_col49[90];
   result_col49[92] <= result_col49[91];
   result_col49[93] <= result_col49[92];
   result_col49[94] <= result_col49[93];
   result_col49[95] <= result_col49[94];
   result_col49[96] <= result_col49[95];
   result_col49[97] <= result_col49[96];
   result_col49[98] <= result_col49[97];
   result_col49[99] <= result_col49[98];
   result_col49[100] <= result_col49[99];
   result_col49[101] <= result_col49[100];
   result_col49[102] <= result_col49[101];
   result_col49[103] <= result_col49[102];
   result_col49[104] <= result_col49[103];
   result_col49[105] <= result_col49[104];
   result_col49[106] <= result_col49[105];
   result_col49[107] <= result_col49[106];
   result_col49[108] <= result_col49[107];
   result_col49[109] <= result_col49[108];
   result_col49[110] <= result_col49[109];
   result_col49[111] <= result_col49[110];
   result_col49[112] <= result_col49[111];
   result_col49[113] <= result_col49[112];
   result_col49[114] <= result_col49[113];
   result_col49[115] <= result_col49[114];
   result_col49[116] <= result_col49[115];
   result_col49[117] <= result_col49[116];

   result_col50[1] <= data_out_4_50;
   result_col50[2] <= result_col50[1];
   result_col50[3] <= result_col50[2];
   result_col50[4] <= result_col50[3];
   result_col50[5] <= result_col50[4];
   result_col50[6] <= result_col50[5];
   result_col50[7] <= result_col50[6];
   result_col50[8] <= result_col50[7];
   result_col50[9] <= result_col50[8];
   result_col50[10] <= result_col50[9];
   result_col50[11] <= result_col50[10];
   result_col50[12] <= result_col50[11];
   result_col50[13] <= result_col50[12];
   result_col50[14] <= result_col50[13];
   result_col50[15] <= result_col50[14];
   result_col50[16] <= result_col50[15];
   result_col50[17] <= result_col50[16];
   result_col50[18] <= result_col50[17];
   result_col50[19] <= result_col50[18];
   result_col50[20] <= result_col50[19];
   result_col50[21] <= result_col50[20];
   result_col50[22] <= result_col50[21];
   result_col50[23] <= result_col50[22];
   result_col50[24] <= result_col50[23];
   result_col50[25] <= result_col50[24];
   result_col50[26] <= result_col50[25];
   result_col50[27] <= result_col50[26];
   result_col50[28] <= result_col50[27];
   result_col50[29] <= result_col50[28];
   result_col50[30] <= result_col50[29];
   result_col50[31] <= result_col50[30];
   result_col50[32] <= result_col50[31];
   result_col50[33] <= result_col50[32];
   result_col50[34] <= result_col50[33];
   result_col50[35] <= result_col50[34];
   result_col50[36] <= result_col50[35];
   result_col50[37] <= result_col50[36];
   result_col50[38] <= result_col50[37];
   result_col50[39] <= result_col50[38];
   result_col50[40] <= result_col50[39];
   result_col50[41] <= result_col50[40];
   result_col50[42] <= result_col50[41];
   result_col50[43] <= result_col50[42];
   result_col50[44] <= result_col50[43];
   result_col50[45] <= result_col50[44];
   result_col50[46] <= result_col50[45];
   result_col50[47] <= result_col50[46];
   result_col50[48] <= result_col50[47];
   result_col50[49] <= result_col50[48];
   result_col50[50] <= result_col50[49];
   result_col50[51] <= result_col50[50];
   result_col50[52] <= result_col50[51];
   result_col50[53] <= result_col50[52];
   result_col50[54] <= result_col50[53];
   result_col50[55] <= result_col50[54];
   result_col50[56] <= result_col50[55];
   result_col50[57] <= result_col50[56];
   result_col50[58] <= result_col50[57];
   result_col50[59] <= result_col50[58];
   result_col50[60] <= result_col50[59];
   result_col50[61] <= result_col50[60];
   result_col50[62] <= result_col50[61];
   result_col50[63] <= result_col50[62];
   result_col50[64] <= result_col50[63];
   result_col50[65] <= result_col50[64];
   result_col50[66] <= result_col50[65];
   result_col50[67] <= result_col50[66];
   result_col50[68] <= result_col50[67];
   result_col50[69] <= result_col50[68];
   result_col50[70] <= result_col50[69];
   result_col50[71] <= result_col50[70];
   result_col50[72] <= result_col50[71];
   result_col50[73] <= result_col50[72];
   result_col50[74] <= result_col50[73];
   result_col50[75] <= result_col50[74];
   result_col50[76] <= result_col50[75];
   result_col50[77] <= result_col50[76];
   result_col50[78] <= result_col50[77];
   result_col50[79] <= result_col50[78];
   result_col50[80] <= result_col50[79];
   result_col50[81] <= result_col50[80];
   result_col50[82] <= result_col50[81];
   result_col50[83] <= result_col50[82];
   result_col50[84] <= result_col50[83];
   result_col50[85] <= result_col50[84];
   result_col50[86] <= result_col50[85];
   result_col50[87] <= result_col50[86];
   result_col50[88] <= result_col50[87];
   result_col50[89] <= result_col50[88];
   result_col50[90] <= result_col50[89];
   result_col50[91] <= result_col50[90];
   result_col50[92] <= result_col50[91];
   result_col50[93] <= result_col50[92];
   result_col50[94] <= result_col50[93];
   result_col50[95] <= result_col50[94];
   result_col50[96] <= result_col50[95];
   result_col50[97] <= result_col50[96];
   result_col50[98] <= result_col50[97];
   result_col50[99] <= result_col50[98];
   result_col50[100] <= result_col50[99];
   result_col50[101] <= result_col50[100];
   result_col50[102] <= result_col50[101];
   result_col50[103] <= result_col50[102];
   result_col50[104] <= result_col50[103];
   result_col50[105] <= result_col50[104];
   result_col50[106] <= result_col50[105];
   result_col50[107] <= result_col50[106];
   result_col50[108] <= result_col50[107];
   result_col50[109] <= result_col50[108];
   result_col50[110] <= result_col50[109];
   result_col50[111] <= result_col50[110];
   result_col50[112] <= result_col50[111];
   result_col50[113] <= result_col50[112];
   result_col50[114] <= result_col50[113];
   result_col50[115] <= result_col50[114];
   result_col50[116] <= result_col50[115];

   result_col51[1] <= data_out_4_51;
   result_col51[2] <= result_col51[1];
   result_col51[3] <= result_col51[2];
   result_col51[4] <= result_col51[3];
   result_col51[5] <= result_col51[4];
   result_col51[6] <= result_col51[5];
   result_col51[7] <= result_col51[6];
   result_col51[8] <= result_col51[7];
   result_col51[9] <= result_col51[8];
   result_col51[10] <= result_col51[9];
   result_col51[11] <= result_col51[10];
   result_col51[12] <= result_col51[11];
   result_col51[13] <= result_col51[12];
   result_col51[14] <= result_col51[13];
   result_col51[15] <= result_col51[14];
   result_col51[16] <= result_col51[15];
   result_col51[17] <= result_col51[16];
   result_col51[18] <= result_col51[17];
   result_col51[19] <= result_col51[18];
   result_col51[20] <= result_col51[19];
   result_col51[21] <= result_col51[20];
   result_col51[22] <= result_col51[21];
   result_col51[23] <= result_col51[22];
   result_col51[24] <= result_col51[23];
   result_col51[25] <= result_col51[24];
   result_col51[26] <= result_col51[25];
   result_col51[27] <= result_col51[26];
   result_col51[28] <= result_col51[27];
   result_col51[29] <= result_col51[28];
   result_col51[30] <= result_col51[29];
   result_col51[31] <= result_col51[30];
   result_col51[32] <= result_col51[31];
   result_col51[33] <= result_col51[32];
   result_col51[34] <= result_col51[33];
   result_col51[35] <= result_col51[34];
   result_col51[36] <= result_col51[35];
   result_col51[37] <= result_col51[36];
   result_col51[38] <= result_col51[37];
   result_col51[39] <= result_col51[38];
   result_col51[40] <= result_col51[39];
   result_col51[41] <= result_col51[40];
   result_col51[42] <= result_col51[41];
   result_col51[43] <= result_col51[42];
   result_col51[44] <= result_col51[43];
   result_col51[45] <= result_col51[44];
   result_col51[46] <= result_col51[45];
   result_col51[47] <= result_col51[46];
   result_col51[48] <= result_col51[47];
   result_col51[49] <= result_col51[48];
   result_col51[50] <= result_col51[49];
   result_col51[51] <= result_col51[50];
   result_col51[52] <= result_col51[51];
   result_col51[53] <= result_col51[52];
   result_col51[54] <= result_col51[53];
   result_col51[55] <= result_col51[54];
   result_col51[56] <= result_col51[55];
   result_col51[57] <= result_col51[56];
   result_col51[58] <= result_col51[57];
   result_col51[59] <= result_col51[58];
   result_col51[60] <= result_col51[59];
   result_col51[61] <= result_col51[60];
   result_col51[62] <= result_col51[61];
   result_col51[63] <= result_col51[62];
   result_col51[64] <= result_col51[63];
   result_col51[65] <= result_col51[64];
   result_col51[66] <= result_col51[65];
   result_col51[67] <= result_col51[66];
   result_col51[68] <= result_col51[67];
   result_col51[69] <= result_col51[68];
   result_col51[70] <= result_col51[69];
   result_col51[71] <= result_col51[70];
   result_col51[72] <= result_col51[71];
   result_col51[73] <= result_col51[72];
   result_col51[74] <= result_col51[73];
   result_col51[75] <= result_col51[74];
   result_col51[76] <= result_col51[75];
   result_col51[77] <= result_col51[76];
   result_col51[78] <= result_col51[77];
   result_col51[79] <= result_col51[78];
   result_col51[80] <= result_col51[79];
   result_col51[81] <= result_col51[80];
   result_col51[82] <= result_col51[81];
   result_col51[83] <= result_col51[82];
   result_col51[84] <= result_col51[83];
   result_col51[85] <= result_col51[84];
   result_col51[86] <= result_col51[85];
   result_col51[87] <= result_col51[86];
   result_col51[88] <= result_col51[87];
   result_col51[89] <= result_col51[88];
   result_col51[90] <= result_col51[89];
   result_col51[91] <= result_col51[90];
   result_col51[92] <= result_col51[91];
   result_col51[93] <= result_col51[92];
   result_col51[94] <= result_col51[93];
   result_col51[95] <= result_col51[94];
   result_col51[96] <= result_col51[95];
   result_col51[97] <= result_col51[96];
   result_col51[98] <= result_col51[97];
   result_col51[99] <= result_col51[98];
   result_col51[100] <= result_col51[99];
   result_col51[101] <= result_col51[100];
   result_col51[102] <= result_col51[101];
   result_col51[103] <= result_col51[102];
   result_col51[104] <= result_col51[103];
   result_col51[105] <= result_col51[104];
   result_col51[106] <= result_col51[105];
   result_col51[107] <= result_col51[106];
   result_col51[108] <= result_col51[107];
   result_col51[109] <= result_col51[108];
   result_col51[110] <= result_col51[109];
   result_col51[111] <= result_col51[110];
   result_col51[112] <= result_col51[111];
   result_col51[113] <= result_col51[112];
   result_col51[114] <= result_col51[113];
   result_col51[115] <= result_col51[114];

   result_col52[1] <= data_out_4_52;
   result_col52[2] <= result_col52[1];
   result_col52[3] <= result_col52[2];
   result_col52[4] <= result_col52[3];
   result_col52[5] <= result_col52[4];
   result_col52[6] <= result_col52[5];
   result_col52[7] <= result_col52[6];
   result_col52[8] <= result_col52[7];
   result_col52[9] <= result_col52[8];
   result_col52[10] <= result_col52[9];
   result_col52[11] <= result_col52[10];
   result_col52[12] <= result_col52[11];
   result_col52[13] <= result_col52[12];
   result_col52[14] <= result_col52[13];
   result_col52[15] <= result_col52[14];
   result_col52[16] <= result_col52[15];
   result_col52[17] <= result_col52[16];
   result_col52[18] <= result_col52[17];
   result_col52[19] <= result_col52[18];
   result_col52[20] <= result_col52[19];
   result_col52[21] <= result_col52[20];
   result_col52[22] <= result_col52[21];
   result_col52[23] <= result_col52[22];
   result_col52[24] <= result_col52[23];
   result_col52[25] <= result_col52[24];
   result_col52[26] <= result_col52[25];
   result_col52[27] <= result_col52[26];
   result_col52[28] <= result_col52[27];
   result_col52[29] <= result_col52[28];
   result_col52[30] <= result_col52[29];
   result_col52[31] <= result_col52[30];
   result_col52[32] <= result_col52[31];
   result_col52[33] <= result_col52[32];
   result_col52[34] <= result_col52[33];
   result_col52[35] <= result_col52[34];
   result_col52[36] <= result_col52[35];
   result_col52[37] <= result_col52[36];
   result_col52[38] <= result_col52[37];
   result_col52[39] <= result_col52[38];
   result_col52[40] <= result_col52[39];
   result_col52[41] <= result_col52[40];
   result_col52[42] <= result_col52[41];
   result_col52[43] <= result_col52[42];
   result_col52[44] <= result_col52[43];
   result_col52[45] <= result_col52[44];
   result_col52[46] <= result_col52[45];
   result_col52[47] <= result_col52[46];
   result_col52[48] <= result_col52[47];
   result_col52[49] <= result_col52[48];
   result_col52[50] <= result_col52[49];
   result_col52[51] <= result_col52[50];
   result_col52[52] <= result_col52[51];
   result_col52[53] <= result_col52[52];
   result_col52[54] <= result_col52[53];
   result_col52[55] <= result_col52[54];
   result_col52[56] <= result_col52[55];
   result_col52[57] <= result_col52[56];
   result_col52[58] <= result_col52[57];
   result_col52[59] <= result_col52[58];
   result_col52[60] <= result_col52[59];
   result_col52[61] <= result_col52[60];
   result_col52[62] <= result_col52[61];
   result_col52[63] <= result_col52[62];
   result_col52[64] <= result_col52[63];
   result_col52[65] <= result_col52[64];
   result_col52[66] <= result_col52[65];
   result_col52[67] <= result_col52[66];
   result_col52[68] <= result_col52[67];
   result_col52[69] <= result_col52[68];
   result_col52[70] <= result_col52[69];
   result_col52[71] <= result_col52[70];
   result_col52[72] <= result_col52[71];
   result_col52[73] <= result_col52[72];
   result_col52[74] <= result_col52[73];
   result_col52[75] <= result_col52[74];
   result_col52[76] <= result_col52[75];
   result_col52[77] <= result_col52[76];
   result_col52[78] <= result_col52[77];
   result_col52[79] <= result_col52[78];
   result_col52[80] <= result_col52[79];
   result_col52[81] <= result_col52[80];
   result_col52[82] <= result_col52[81];
   result_col52[83] <= result_col52[82];
   result_col52[84] <= result_col52[83];
   result_col52[85] <= result_col52[84];
   result_col52[86] <= result_col52[85];
   result_col52[87] <= result_col52[86];
   result_col52[88] <= result_col52[87];
   result_col52[89] <= result_col52[88];
   result_col52[90] <= result_col52[89];
   result_col52[91] <= result_col52[90];
   result_col52[92] <= result_col52[91];
   result_col52[93] <= result_col52[92];
   result_col52[94] <= result_col52[93];
   result_col52[95] <= result_col52[94];
   result_col52[96] <= result_col52[95];
   result_col52[97] <= result_col52[96];
   result_col52[98] <= result_col52[97];
   result_col52[99] <= result_col52[98];
   result_col52[100] <= result_col52[99];
   result_col52[101] <= result_col52[100];
   result_col52[102] <= result_col52[101];
   result_col52[103] <= result_col52[102];
   result_col52[104] <= result_col52[103];
   result_col52[105] <= result_col52[104];
   result_col52[106] <= result_col52[105];
   result_col52[107] <= result_col52[106];
   result_col52[108] <= result_col52[107];
   result_col52[109] <= result_col52[108];
   result_col52[110] <= result_col52[109];
   result_col52[111] <= result_col52[110];
   result_col52[112] <= result_col52[111];
   result_col52[113] <= result_col52[112];
   result_col52[114] <= result_col52[113];

   result_col53[1] <= data_out_4_53;
   result_col53[2] <= result_col53[1];
   result_col53[3] <= result_col53[2];
   result_col53[4] <= result_col53[3];
   result_col53[5] <= result_col53[4];
   result_col53[6] <= result_col53[5];
   result_col53[7] <= result_col53[6];
   result_col53[8] <= result_col53[7];
   result_col53[9] <= result_col53[8];
   result_col53[10] <= result_col53[9];
   result_col53[11] <= result_col53[10];
   result_col53[12] <= result_col53[11];
   result_col53[13] <= result_col53[12];
   result_col53[14] <= result_col53[13];
   result_col53[15] <= result_col53[14];
   result_col53[16] <= result_col53[15];
   result_col53[17] <= result_col53[16];
   result_col53[18] <= result_col53[17];
   result_col53[19] <= result_col53[18];
   result_col53[20] <= result_col53[19];
   result_col53[21] <= result_col53[20];
   result_col53[22] <= result_col53[21];
   result_col53[23] <= result_col53[22];
   result_col53[24] <= result_col53[23];
   result_col53[25] <= result_col53[24];
   result_col53[26] <= result_col53[25];
   result_col53[27] <= result_col53[26];
   result_col53[28] <= result_col53[27];
   result_col53[29] <= result_col53[28];
   result_col53[30] <= result_col53[29];
   result_col53[31] <= result_col53[30];
   result_col53[32] <= result_col53[31];
   result_col53[33] <= result_col53[32];
   result_col53[34] <= result_col53[33];
   result_col53[35] <= result_col53[34];
   result_col53[36] <= result_col53[35];
   result_col53[37] <= result_col53[36];
   result_col53[38] <= result_col53[37];
   result_col53[39] <= result_col53[38];
   result_col53[40] <= result_col53[39];
   result_col53[41] <= result_col53[40];
   result_col53[42] <= result_col53[41];
   result_col53[43] <= result_col53[42];
   result_col53[44] <= result_col53[43];
   result_col53[45] <= result_col53[44];
   result_col53[46] <= result_col53[45];
   result_col53[47] <= result_col53[46];
   result_col53[48] <= result_col53[47];
   result_col53[49] <= result_col53[48];
   result_col53[50] <= result_col53[49];
   result_col53[51] <= result_col53[50];
   result_col53[52] <= result_col53[51];
   result_col53[53] <= result_col53[52];
   result_col53[54] <= result_col53[53];
   result_col53[55] <= result_col53[54];
   result_col53[56] <= result_col53[55];
   result_col53[57] <= result_col53[56];
   result_col53[58] <= result_col53[57];
   result_col53[59] <= result_col53[58];
   result_col53[60] <= result_col53[59];
   result_col53[61] <= result_col53[60];
   result_col53[62] <= result_col53[61];
   result_col53[63] <= result_col53[62];
   result_col53[64] <= result_col53[63];
   result_col53[65] <= result_col53[64];
   result_col53[66] <= result_col53[65];
   result_col53[67] <= result_col53[66];
   result_col53[68] <= result_col53[67];
   result_col53[69] <= result_col53[68];
   result_col53[70] <= result_col53[69];
   result_col53[71] <= result_col53[70];
   result_col53[72] <= result_col53[71];
   result_col53[73] <= result_col53[72];
   result_col53[74] <= result_col53[73];
   result_col53[75] <= result_col53[74];
   result_col53[76] <= result_col53[75];
   result_col53[77] <= result_col53[76];
   result_col53[78] <= result_col53[77];
   result_col53[79] <= result_col53[78];
   result_col53[80] <= result_col53[79];
   result_col53[81] <= result_col53[80];
   result_col53[82] <= result_col53[81];
   result_col53[83] <= result_col53[82];
   result_col53[84] <= result_col53[83];
   result_col53[85] <= result_col53[84];
   result_col53[86] <= result_col53[85];
   result_col53[87] <= result_col53[86];
   result_col53[88] <= result_col53[87];
   result_col53[89] <= result_col53[88];
   result_col53[90] <= result_col53[89];
   result_col53[91] <= result_col53[90];
   result_col53[92] <= result_col53[91];
   result_col53[93] <= result_col53[92];
   result_col53[94] <= result_col53[93];
   result_col53[95] <= result_col53[94];
   result_col53[96] <= result_col53[95];
   result_col53[97] <= result_col53[96];
   result_col53[98] <= result_col53[97];
   result_col53[99] <= result_col53[98];
   result_col53[100] <= result_col53[99];
   result_col53[101] <= result_col53[100];
   result_col53[102] <= result_col53[101];
   result_col53[103] <= result_col53[102];
   result_col53[104] <= result_col53[103];
   result_col53[105] <= result_col53[104];
   result_col53[106] <= result_col53[105];
   result_col53[107] <= result_col53[106];
   result_col53[108] <= result_col53[107];
   result_col53[109] <= result_col53[108];
   result_col53[110] <= result_col53[109];
   result_col53[111] <= result_col53[110];
   result_col53[112] <= result_col53[111];
   result_col53[113] <= result_col53[112];

   result_col54[1] <= data_out_4_54;
   result_col54[2] <= result_col54[1];
   result_col54[3] <= result_col54[2];
   result_col54[4] <= result_col54[3];
   result_col54[5] <= result_col54[4];
   result_col54[6] <= result_col54[5];
   result_col54[7] <= result_col54[6];
   result_col54[8] <= result_col54[7];
   result_col54[9] <= result_col54[8];
   result_col54[10] <= result_col54[9];
   result_col54[11] <= result_col54[10];
   result_col54[12] <= result_col54[11];
   result_col54[13] <= result_col54[12];
   result_col54[14] <= result_col54[13];
   result_col54[15] <= result_col54[14];
   result_col54[16] <= result_col54[15];
   result_col54[17] <= result_col54[16];
   result_col54[18] <= result_col54[17];
   result_col54[19] <= result_col54[18];
   result_col54[20] <= result_col54[19];
   result_col54[21] <= result_col54[20];
   result_col54[22] <= result_col54[21];
   result_col54[23] <= result_col54[22];
   result_col54[24] <= result_col54[23];
   result_col54[25] <= result_col54[24];
   result_col54[26] <= result_col54[25];
   result_col54[27] <= result_col54[26];
   result_col54[28] <= result_col54[27];
   result_col54[29] <= result_col54[28];
   result_col54[30] <= result_col54[29];
   result_col54[31] <= result_col54[30];
   result_col54[32] <= result_col54[31];
   result_col54[33] <= result_col54[32];
   result_col54[34] <= result_col54[33];
   result_col54[35] <= result_col54[34];
   result_col54[36] <= result_col54[35];
   result_col54[37] <= result_col54[36];
   result_col54[38] <= result_col54[37];
   result_col54[39] <= result_col54[38];
   result_col54[40] <= result_col54[39];
   result_col54[41] <= result_col54[40];
   result_col54[42] <= result_col54[41];
   result_col54[43] <= result_col54[42];
   result_col54[44] <= result_col54[43];
   result_col54[45] <= result_col54[44];
   result_col54[46] <= result_col54[45];
   result_col54[47] <= result_col54[46];
   result_col54[48] <= result_col54[47];
   result_col54[49] <= result_col54[48];
   result_col54[50] <= result_col54[49];
   result_col54[51] <= result_col54[50];
   result_col54[52] <= result_col54[51];
   result_col54[53] <= result_col54[52];
   result_col54[54] <= result_col54[53];
   result_col54[55] <= result_col54[54];
   result_col54[56] <= result_col54[55];
   result_col54[57] <= result_col54[56];
   result_col54[58] <= result_col54[57];
   result_col54[59] <= result_col54[58];
   result_col54[60] <= result_col54[59];
   result_col54[61] <= result_col54[60];
   result_col54[62] <= result_col54[61];
   result_col54[63] <= result_col54[62];
   result_col54[64] <= result_col54[63];
   result_col54[65] <= result_col54[64];
   result_col54[66] <= result_col54[65];
   result_col54[67] <= result_col54[66];
   result_col54[68] <= result_col54[67];
   result_col54[69] <= result_col54[68];
   result_col54[70] <= result_col54[69];
   result_col54[71] <= result_col54[70];
   result_col54[72] <= result_col54[71];
   result_col54[73] <= result_col54[72];
   result_col54[74] <= result_col54[73];
   result_col54[75] <= result_col54[74];
   result_col54[76] <= result_col54[75];
   result_col54[77] <= result_col54[76];
   result_col54[78] <= result_col54[77];
   result_col54[79] <= result_col54[78];
   result_col54[80] <= result_col54[79];
   result_col54[81] <= result_col54[80];
   result_col54[82] <= result_col54[81];
   result_col54[83] <= result_col54[82];
   result_col54[84] <= result_col54[83];
   result_col54[85] <= result_col54[84];
   result_col54[86] <= result_col54[85];
   result_col54[87] <= result_col54[86];
   result_col54[88] <= result_col54[87];
   result_col54[89] <= result_col54[88];
   result_col54[90] <= result_col54[89];
   result_col54[91] <= result_col54[90];
   result_col54[92] <= result_col54[91];
   result_col54[93] <= result_col54[92];
   result_col54[94] <= result_col54[93];
   result_col54[95] <= result_col54[94];
   result_col54[96] <= result_col54[95];
   result_col54[97] <= result_col54[96];
   result_col54[98] <= result_col54[97];
   result_col54[99] <= result_col54[98];
   result_col54[100] <= result_col54[99];
   result_col54[101] <= result_col54[100];
   result_col54[102] <= result_col54[101];
   result_col54[103] <= result_col54[102];
   result_col54[104] <= result_col54[103];
   result_col54[105] <= result_col54[104];
   result_col54[106] <= result_col54[105];
   result_col54[107] <= result_col54[106];
   result_col54[108] <= result_col54[107];
   result_col54[109] <= result_col54[108];
   result_col54[110] <= result_col54[109];
   result_col54[111] <= result_col54[110];
   result_col54[112] <= result_col54[111];

   result_col55[1] <= data_out_4_55;
   result_col55[2] <= result_col55[1];
   result_col55[3] <= result_col55[2];
   result_col55[4] <= result_col55[3];
   result_col55[5] <= result_col55[4];
   result_col55[6] <= result_col55[5];
   result_col55[7] <= result_col55[6];
   result_col55[8] <= result_col55[7];
   result_col55[9] <= result_col55[8];
   result_col55[10] <= result_col55[9];
   result_col55[11] <= result_col55[10];
   result_col55[12] <= result_col55[11];
   result_col55[13] <= result_col55[12];
   result_col55[14] <= result_col55[13];
   result_col55[15] <= result_col55[14];
   result_col55[16] <= result_col55[15];
   result_col55[17] <= result_col55[16];
   result_col55[18] <= result_col55[17];
   result_col55[19] <= result_col55[18];
   result_col55[20] <= result_col55[19];
   result_col55[21] <= result_col55[20];
   result_col55[22] <= result_col55[21];
   result_col55[23] <= result_col55[22];
   result_col55[24] <= result_col55[23];
   result_col55[25] <= result_col55[24];
   result_col55[26] <= result_col55[25];
   result_col55[27] <= result_col55[26];
   result_col55[28] <= result_col55[27];
   result_col55[29] <= result_col55[28];
   result_col55[30] <= result_col55[29];
   result_col55[31] <= result_col55[30];
   result_col55[32] <= result_col55[31];
   result_col55[33] <= result_col55[32];
   result_col55[34] <= result_col55[33];
   result_col55[35] <= result_col55[34];
   result_col55[36] <= result_col55[35];
   result_col55[37] <= result_col55[36];
   result_col55[38] <= result_col55[37];
   result_col55[39] <= result_col55[38];
   result_col55[40] <= result_col55[39];
   result_col55[41] <= result_col55[40];
   result_col55[42] <= result_col55[41];
   result_col55[43] <= result_col55[42];
   result_col55[44] <= result_col55[43];
   result_col55[45] <= result_col55[44];
   result_col55[46] <= result_col55[45];
   result_col55[47] <= result_col55[46];
   result_col55[48] <= result_col55[47];
   result_col55[49] <= result_col55[48];
   result_col55[50] <= result_col55[49];
   result_col55[51] <= result_col55[50];
   result_col55[52] <= result_col55[51];
   result_col55[53] <= result_col55[52];
   result_col55[54] <= result_col55[53];
   result_col55[55] <= result_col55[54];
   result_col55[56] <= result_col55[55];
   result_col55[57] <= result_col55[56];
   result_col55[58] <= result_col55[57];
   result_col55[59] <= result_col55[58];
   result_col55[60] <= result_col55[59];
   result_col55[61] <= result_col55[60];
   result_col55[62] <= result_col55[61];
   result_col55[63] <= result_col55[62];
   result_col55[64] <= result_col55[63];
   result_col55[65] <= result_col55[64];
   result_col55[66] <= result_col55[65];
   result_col55[67] <= result_col55[66];
   result_col55[68] <= result_col55[67];
   result_col55[69] <= result_col55[68];
   result_col55[70] <= result_col55[69];
   result_col55[71] <= result_col55[70];
   result_col55[72] <= result_col55[71];
   result_col55[73] <= result_col55[72];
   result_col55[74] <= result_col55[73];
   result_col55[75] <= result_col55[74];
   result_col55[76] <= result_col55[75];
   result_col55[77] <= result_col55[76];
   result_col55[78] <= result_col55[77];
   result_col55[79] <= result_col55[78];
   result_col55[80] <= result_col55[79];
   result_col55[81] <= result_col55[80];
   result_col55[82] <= result_col55[81];
   result_col55[83] <= result_col55[82];
   result_col55[84] <= result_col55[83];
   result_col55[85] <= result_col55[84];
   result_col55[86] <= result_col55[85];
   result_col55[87] <= result_col55[86];
   result_col55[88] <= result_col55[87];
   result_col55[89] <= result_col55[88];
   result_col55[90] <= result_col55[89];
   result_col55[91] <= result_col55[90];
   result_col55[92] <= result_col55[91];
   result_col55[93] <= result_col55[92];
   result_col55[94] <= result_col55[93];
   result_col55[95] <= result_col55[94];
   result_col55[96] <= result_col55[95];
   result_col55[97] <= result_col55[96];
   result_col55[98] <= result_col55[97];
   result_col55[99] <= result_col55[98];
   result_col55[100] <= result_col55[99];
   result_col55[101] <= result_col55[100];
   result_col55[102] <= result_col55[101];
   result_col55[103] <= result_col55[102];
   result_col55[104] <= result_col55[103];
   result_col55[105] <= result_col55[104];
   result_col55[106] <= result_col55[105];
   result_col55[107] <= result_col55[106];
   result_col55[108] <= result_col55[107];
   result_col55[109] <= result_col55[108];
   result_col55[110] <= result_col55[109];
   result_col55[111] <= result_col55[110];

   result_col56[1] <= data_out_4_56;
   result_col56[2] <= result_col56[1];
   result_col56[3] <= result_col56[2];
   result_col56[4] <= result_col56[3];
   result_col56[5] <= result_col56[4];
   result_col56[6] <= result_col56[5];
   result_col56[7] <= result_col56[6];
   result_col56[8] <= result_col56[7];
   result_col56[9] <= result_col56[8];
   result_col56[10] <= result_col56[9];
   result_col56[11] <= result_col56[10];
   result_col56[12] <= result_col56[11];
   result_col56[13] <= result_col56[12];
   result_col56[14] <= result_col56[13];
   result_col56[15] <= result_col56[14];
   result_col56[16] <= result_col56[15];
   result_col56[17] <= result_col56[16];
   result_col56[18] <= result_col56[17];
   result_col56[19] <= result_col56[18];
   result_col56[20] <= result_col56[19];
   result_col56[21] <= result_col56[20];
   result_col56[22] <= result_col56[21];
   result_col56[23] <= result_col56[22];
   result_col56[24] <= result_col56[23];
   result_col56[25] <= result_col56[24];
   result_col56[26] <= result_col56[25];
   result_col56[27] <= result_col56[26];
   result_col56[28] <= result_col56[27];
   result_col56[29] <= result_col56[28];
   result_col56[30] <= result_col56[29];
   result_col56[31] <= result_col56[30];
   result_col56[32] <= result_col56[31];
   result_col56[33] <= result_col56[32];
   result_col56[34] <= result_col56[33];
   result_col56[35] <= result_col56[34];
   result_col56[36] <= result_col56[35];
   result_col56[37] <= result_col56[36];
   result_col56[38] <= result_col56[37];
   result_col56[39] <= result_col56[38];
   result_col56[40] <= result_col56[39];
   result_col56[41] <= result_col56[40];
   result_col56[42] <= result_col56[41];
   result_col56[43] <= result_col56[42];
   result_col56[44] <= result_col56[43];
   result_col56[45] <= result_col56[44];
   result_col56[46] <= result_col56[45];
   result_col56[47] <= result_col56[46];
   result_col56[48] <= result_col56[47];
   result_col56[49] <= result_col56[48];
   result_col56[50] <= result_col56[49];
   result_col56[51] <= result_col56[50];
   result_col56[52] <= result_col56[51];
   result_col56[53] <= result_col56[52];
   result_col56[54] <= result_col56[53];
   result_col56[55] <= result_col56[54];
   result_col56[56] <= result_col56[55];
   result_col56[57] <= result_col56[56];
   result_col56[58] <= result_col56[57];
   result_col56[59] <= result_col56[58];
   result_col56[60] <= result_col56[59];
   result_col56[61] <= result_col56[60];
   result_col56[62] <= result_col56[61];
   result_col56[63] <= result_col56[62];
   result_col56[64] <= result_col56[63];
   result_col56[65] <= result_col56[64];
   result_col56[66] <= result_col56[65];
   result_col56[67] <= result_col56[66];
   result_col56[68] <= result_col56[67];
   result_col56[69] <= result_col56[68];
   result_col56[70] <= result_col56[69];
   result_col56[71] <= result_col56[70];
   result_col56[72] <= result_col56[71];
   result_col56[73] <= result_col56[72];
   result_col56[74] <= result_col56[73];
   result_col56[75] <= result_col56[74];
   result_col56[76] <= result_col56[75];
   result_col56[77] <= result_col56[76];
   result_col56[78] <= result_col56[77];
   result_col56[79] <= result_col56[78];
   result_col56[80] <= result_col56[79];
   result_col56[81] <= result_col56[80];
   result_col56[82] <= result_col56[81];
   result_col56[83] <= result_col56[82];
   result_col56[84] <= result_col56[83];
   result_col56[85] <= result_col56[84];
   result_col56[86] <= result_col56[85];
   result_col56[87] <= result_col56[86];
   result_col56[88] <= result_col56[87];
   result_col56[89] <= result_col56[88];
   result_col56[90] <= result_col56[89];
   result_col56[91] <= result_col56[90];
   result_col56[92] <= result_col56[91];
   result_col56[93] <= result_col56[92];
   result_col56[94] <= result_col56[93];
   result_col56[95] <= result_col56[94];
   result_col56[96] <= result_col56[95];
   result_col56[97] <= result_col56[96];
   result_col56[98] <= result_col56[97];
   result_col56[99] <= result_col56[98];
   result_col56[100] <= result_col56[99];
   result_col56[101] <= result_col56[100];
   result_col56[102] <= result_col56[101];
   result_col56[103] <= result_col56[102];
   result_col56[104] <= result_col56[103];
   result_col56[105] <= result_col56[104];
   result_col56[106] <= result_col56[105];
   result_col56[107] <= result_col56[106];
   result_col56[108] <= result_col56[107];
   result_col56[109] <= result_col56[108];
   result_col56[110] <= result_col56[109];

   result_col57[1] <= data_out_4_57;
   result_col57[2] <= result_col57[1];
   result_col57[3] <= result_col57[2];
   result_col57[4] <= result_col57[3];
   result_col57[5] <= result_col57[4];
   result_col57[6] <= result_col57[5];
   result_col57[7] <= result_col57[6];
   result_col57[8] <= result_col57[7];
   result_col57[9] <= result_col57[8];
   result_col57[10] <= result_col57[9];
   result_col57[11] <= result_col57[10];
   result_col57[12] <= result_col57[11];
   result_col57[13] <= result_col57[12];
   result_col57[14] <= result_col57[13];
   result_col57[15] <= result_col57[14];
   result_col57[16] <= result_col57[15];
   result_col57[17] <= result_col57[16];
   result_col57[18] <= result_col57[17];
   result_col57[19] <= result_col57[18];
   result_col57[20] <= result_col57[19];
   result_col57[21] <= result_col57[20];
   result_col57[22] <= result_col57[21];
   result_col57[23] <= result_col57[22];
   result_col57[24] <= result_col57[23];
   result_col57[25] <= result_col57[24];
   result_col57[26] <= result_col57[25];
   result_col57[27] <= result_col57[26];
   result_col57[28] <= result_col57[27];
   result_col57[29] <= result_col57[28];
   result_col57[30] <= result_col57[29];
   result_col57[31] <= result_col57[30];
   result_col57[32] <= result_col57[31];
   result_col57[33] <= result_col57[32];
   result_col57[34] <= result_col57[33];
   result_col57[35] <= result_col57[34];
   result_col57[36] <= result_col57[35];
   result_col57[37] <= result_col57[36];
   result_col57[38] <= result_col57[37];
   result_col57[39] <= result_col57[38];
   result_col57[40] <= result_col57[39];
   result_col57[41] <= result_col57[40];
   result_col57[42] <= result_col57[41];
   result_col57[43] <= result_col57[42];
   result_col57[44] <= result_col57[43];
   result_col57[45] <= result_col57[44];
   result_col57[46] <= result_col57[45];
   result_col57[47] <= result_col57[46];
   result_col57[48] <= result_col57[47];
   result_col57[49] <= result_col57[48];
   result_col57[50] <= result_col57[49];
   result_col57[51] <= result_col57[50];
   result_col57[52] <= result_col57[51];
   result_col57[53] <= result_col57[52];
   result_col57[54] <= result_col57[53];
   result_col57[55] <= result_col57[54];
   result_col57[56] <= result_col57[55];
   result_col57[57] <= result_col57[56];
   result_col57[58] <= result_col57[57];
   result_col57[59] <= result_col57[58];
   result_col57[60] <= result_col57[59];
   result_col57[61] <= result_col57[60];
   result_col57[62] <= result_col57[61];
   result_col57[63] <= result_col57[62];
   result_col57[64] <= result_col57[63];
   result_col57[65] <= result_col57[64];
   result_col57[66] <= result_col57[65];
   result_col57[67] <= result_col57[66];
   result_col57[68] <= result_col57[67];
   result_col57[69] <= result_col57[68];
   result_col57[70] <= result_col57[69];
   result_col57[71] <= result_col57[70];
   result_col57[72] <= result_col57[71];
   result_col57[73] <= result_col57[72];
   result_col57[74] <= result_col57[73];
   result_col57[75] <= result_col57[74];
   result_col57[76] <= result_col57[75];
   result_col57[77] <= result_col57[76];
   result_col57[78] <= result_col57[77];
   result_col57[79] <= result_col57[78];
   result_col57[80] <= result_col57[79];
   result_col57[81] <= result_col57[80];
   result_col57[82] <= result_col57[81];
   result_col57[83] <= result_col57[82];
   result_col57[84] <= result_col57[83];
   result_col57[85] <= result_col57[84];
   result_col57[86] <= result_col57[85];
   result_col57[87] <= result_col57[86];
   result_col57[88] <= result_col57[87];
   result_col57[89] <= result_col57[88];
   result_col57[90] <= result_col57[89];
   result_col57[91] <= result_col57[90];
   result_col57[92] <= result_col57[91];
   result_col57[93] <= result_col57[92];
   result_col57[94] <= result_col57[93];
   result_col57[95] <= result_col57[94];
   result_col57[96] <= result_col57[95];
   result_col57[97] <= result_col57[96];
   result_col57[98] <= result_col57[97];
   result_col57[99] <= result_col57[98];
   result_col57[100] <= result_col57[99];
   result_col57[101] <= result_col57[100];
   result_col57[102] <= result_col57[101];
   result_col57[103] <= result_col57[102];
   result_col57[104] <= result_col57[103];
   result_col57[105] <= result_col57[104];
   result_col57[106] <= result_col57[105];
   result_col57[107] <= result_col57[106];
   result_col57[108] <= result_col57[107];
   result_col57[109] <= result_col57[108];

   result_col58[1] <= data_out_4_58;
   result_col58[2] <= result_col58[1];
   result_col58[3] <= result_col58[2];
   result_col58[4] <= result_col58[3];
   result_col58[5] <= result_col58[4];
   result_col58[6] <= result_col58[5];
   result_col58[7] <= result_col58[6];
   result_col58[8] <= result_col58[7];
   result_col58[9] <= result_col58[8];
   result_col58[10] <= result_col58[9];
   result_col58[11] <= result_col58[10];
   result_col58[12] <= result_col58[11];
   result_col58[13] <= result_col58[12];
   result_col58[14] <= result_col58[13];
   result_col58[15] <= result_col58[14];
   result_col58[16] <= result_col58[15];
   result_col58[17] <= result_col58[16];
   result_col58[18] <= result_col58[17];
   result_col58[19] <= result_col58[18];
   result_col58[20] <= result_col58[19];
   result_col58[21] <= result_col58[20];
   result_col58[22] <= result_col58[21];
   result_col58[23] <= result_col58[22];
   result_col58[24] <= result_col58[23];
   result_col58[25] <= result_col58[24];
   result_col58[26] <= result_col58[25];
   result_col58[27] <= result_col58[26];
   result_col58[28] <= result_col58[27];
   result_col58[29] <= result_col58[28];
   result_col58[30] <= result_col58[29];
   result_col58[31] <= result_col58[30];
   result_col58[32] <= result_col58[31];
   result_col58[33] <= result_col58[32];
   result_col58[34] <= result_col58[33];
   result_col58[35] <= result_col58[34];
   result_col58[36] <= result_col58[35];
   result_col58[37] <= result_col58[36];
   result_col58[38] <= result_col58[37];
   result_col58[39] <= result_col58[38];
   result_col58[40] <= result_col58[39];
   result_col58[41] <= result_col58[40];
   result_col58[42] <= result_col58[41];
   result_col58[43] <= result_col58[42];
   result_col58[44] <= result_col58[43];
   result_col58[45] <= result_col58[44];
   result_col58[46] <= result_col58[45];
   result_col58[47] <= result_col58[46];
   result_col58[48] <= result_col58[47];
   result_col58[49] <= result_col58[48];
   result_col58[50] <= result_col58[49];
   result_col58[51] <= result_col58[50];
   result_col58[52] <= result_col58[51];
   result_col58[53] <= result_col58[52];
   result_col58[54] <= result_col58[53];
   result_col58[55] <= result_col58[54];
   result_col58[56] <= result_col58[55];
   result_col58[57] <= result_col58[56];
   result_col58[58] <= result_col58[57];
   result_col58[59] <= result_col58[58];
   result_col58[60] <= result_col58[59];
   result_col58[61] <= result_col58[60];
   result_col58[62] <= result_col58[61];
   result_col58[63] <= result_col58[62];
   result_col58[64] <= result_col58[63];
   result_col58[65] <= result_col58[64];
   result_col58[66] <= result_col58[65];
   result_col58[67] <= result_col58[66];
   result_col58[68] <= result_col58[67];
   result_col58[69] <= result_col58[68];
   result_col58[70] <= result_col58[69];
   result_col58[71] <= result_col58[70];
   result_col58[72] <= result_col58[71];
   result_col58[73] <= result_col58[72];
   result_col58[74] <= result_col58[73];
   result_col58[75] <= result_col58[74];
   result_col58[76] <= result_col58[75];
   result_col58[77] <= result_col58[76];
   result_col58[78] <= result_col58[77];
   result_col58[79] <= result_col58[78];
   result_col58[80] <= result_col58[79];
   result_col58[81] <= result_col58[80];
   result_col58[82] <= result_col58[81];
   result_col58[83] <= result_col58[82];
   result_col58[84] <= result_col58[83];
   result_col58[85] <= result_col58[84];
   result_col58[86] <= result_col58[85];
   result_col58[87] <= result_col58[86];
   result_col58[88] <= result_col58[87];
   result_col58[89] <= result_col58[88];
   result_col58[90] <= result_col58[89];
   result_col58[91] <= result_col58[90];
   result_col58[92] <= result_col58[91];
   result_col58[93] <= result_col58[92];
   result_col58[94] <= result_col58[93];
   result_col58[95] <= result_col58[94];
   result_col58[96] <= result_col58[95];
   result_col58[97] <= result_col58[96];
   result_col58[98] <= result_col58[97];
   result_col58[99] <= result_col58[98];
   result_col58[100] <= result_col58[99];
   result_col58[101] <= result_col58[100];
   result_col58[102] <= result_col58[101];
   result_col58[103] <= result_col58[102];
   result_col58[104] <= result_col58[103];
   result_col58[105] <= result_col58[104];
   result_col58[106] <= result_col58[105];
   result_col58[107] <= result_col58[106];
   result_col58[108] <= result_col58[107];

   result_col59[1] <= data_out_4_59;
   result_col59[2] <= result_col59[1];
   result_col59[3] <= result_col59[2];
   result_col59[4] <= result_col59[3];
   result_col59[5] <= result_col59[4];
   result_col59[6] <= result_col59[5];
   result_col59[7] <= result_col59[6];
   result_col59[8] <= result_col59[7];
   result_col59[9] <= result_col59[8];
   result_col59[10] <= result_col59[9];
   result_col59[11] <= result_col59[10];
   result_col59[12] <= result_col59[11];
   result_col59[13] <= result_col59[12];
   result_col59[14] <= result_col59[13];
   result_col59[15] <= result_col59[14];
   result_col59[16] <= result_col59[15];
   result_col59[17] <= result_col59[16];
   result_col59[18] <= result_col59[17];
   result_col59[19] <= result_col59[18];
   result_col59[20] <= result_col59[19];
   result_col59[21] <= result_col59[20];
   result_col59[22] <= result_col59[21];
   result_col59[23] <= result_col59[22];
   result_col59[24] <= result_col59[23];
   result_col59[25] <= result_col59[24];
   result_col59[26] <= result_col59[25];
   result_col59[27] <= result_col59[26];
   result_col59[28] <= result_col59[27];
   result_col59[29] <= result_col59[28];
   result_col59[30] <= result_col59[29];
   result_col59[31] <= result_col59[30];
   result_col59[32] <= result_col59[31];
   result_col59[33] <= result_col59[32];
   result_col59[34] <= result_col59[33];
   result_col59[35] <= result_col59[34];
   result_col59[36] <= result_col59[35];
   result_col59[37] <= result_col59[36];
   result_col59[38] <= result_col59[37];
   result_col59[39] <= result_col59[38];
   result_col59[40] <= result_col59[39];
   result_col59[41] <= result_col59[40];
   result_col59[42] <= result_col59[41];
   result_col59[43] <= result_col59[42];
   result_col59[44] <= result_col59[43];
   result_col59[45] <= result_col59[44];
   result_col59[46] <= result_col59[45];
   result_col59[47] <= result_col59[46];
   result_col59[48] <= result_col59[47];
   result_col59[49] <= result_col59[48];
   result_col59[50] <= result_col59[49];
   result_col59[51] <= result_col59[50];
   result_col59[52] <= result_col59[51];
   result_col59[53] <= result_col59[52];
   result_col59[54] <= result_col59[53];
   result_col59[55] <= result_col59[54];
   result_col59[56] <= result_col59[55];
   result_col59[57] <= result_col59[56];
   result_col59[58] <= result_col59[57];
   result_col59[59] <= result_col59[58];
   result_col59[60] <= result_col59[59];
   result_col59[61] <= result_col59[60];
   result_col59[62] <= result_col59[61];
   result_col59[63] <= result_col59[62];
   result_col59[64] <= result_col59[63];
   result_col59[65] <= result_col59[64];
   result_col59[66] <= result_col59[65];
   result_col59[67] <= result_col59[66];
   result_col59[68] <= result_col59[67];
   result_col59[69] <= result_col59[68];
   result_col59[70] <= result_col59[69];
   result_col59[71] <= result_col59[70];
   result_col59[72] <= result_col59[71];
   result_col59[73] <= result_col59[72];
   result_col59[74] <= result_col59[73];
   result_col59[75] <= result_col59[74];
   result_col59[76] <= result_col59[75];
   result_col59[77] <= result_col59[76];
   result_col59[78] <= result_col59[77];
   result_col59[79] <= result_col59[78];
   result_col59[80] <= result_col59[79];
   result_col59[81] <= result_col59[80];
   result_col59[82] <= result_col59[81];
   result_col59[83] <= result_col59[82];
   result_col59[84] <= result_col59[83];
   result_col59[85] <= result_col59[84];
   result_col59[86] <= result_col59[85];
   result_col59[87] <= result_col59[86];
   result_col59[88] <= result_col59[87];
   result_col59[89] <= result_col59[88];
   result_col59[90] <= result_col59[89];
   result_col59[91] <= result_col59[90];
   result_col59[92] <= result_col59[91];
   result_col59[93] <= result_col59[92];
   result_col59[94] <= result_col59[93];
   result_col59[95] <= result_col59[94];
   result_col59[96] <= result_col59[95];
   result_col59[97] <= result_col59[96];
   result_col59[98] <= result_col59[97];
   result_col59[99] <= result_col59[98];
   result_col59[100] <= result_col59[99];
   result_col59[101] <= result_col59[100];
   result_col59[102] <= result_col59[101];
   result_col59[103] <= result_col59[102];
   result_col59[104] <= result_col59[103];
   result_col59[105] <= result_col59[104];
   result_col59[106] <= result_col59[105];
   result_col59[107] <= result_col59[106];

   result_col60[1] <= data_out_4_60;
   result_col60[2] <= result_col60[1];
   result_col60[3] <= result_col60[2];
   result_col60[4] <= result_col60[3];
   result_col60[5] <= result_col60[4];
   result_col60[6] <= result_col60[5];
   result_col60[7] <= result_col60[6];
   result_col60[8] <= result_col60[7];
   result_col60[9] <= result_col60[8];
   result_col60[10] <= result_col60[9];
   result_col60[11] <= result_col60[10];
   result_col60[12] <= result_col60[11];
   result_col60[13] <= result_col60[12];
   result_col60[14] <= result_col60[13];
   result_col60[15] <= result_col60[14];
   result_col60[16] <= result_col60[15];
   result_col60[17] <= result_col60[16];
   result_col60[18] <= result_col60[17];
   result_col60[19] <= result_col60[18];
   result_col60[20] <= result_col60[19];
   result_col60[21] <= result_col60[20];
   result_col60[22] <= result_col60[21];
   result_col60[23] <= result_col60[22];
   result_col60[24] <= result_col60[23];
   result_col60[25] <= result_col60[24];
   result_col60[26] <= result_col60[25];
   result_col60[27] <= result_col60[26];
   result_col60[28] <= result_col60[27];
   result_col60[29] <= result_col60[28];
   result_col60[30] <= result_col60[29];
   result_col60[31] <= result_col60[30];
   result_col60[32] <= result_col60[31];
   result_col60[33] <= result_col60[32];
   result_col60[34] <= result_col60[33];
   result_col60[35] <= result_col60[34];
   result_col60[36] <= result_col60[35];
   result_col60[37] <= result_col60[36];
   result_col60[38] <= result_col60[37];
   result_col60[39] <= result_col60[38];
   result_col60[40] <= result_col60[39];
   result_col60[41] <= result_col60[40];
   result_col60[42] <= result_col60[41];
   result_col60[43] <= result_col60[42];
   result_col60[44] <= result_col60[43];
   result_col60[45] <= result_col60[44];
   result_col60[46] <= result_col60[45];
   result_col60[47] <= result_col60[46];
   result_col60[48] <= result_col60[47];
   result_col60[49] <= result_col60[48];
   result_col60[50] <= result_col60[49];
   result_col60[51] <= result_col60[50];
   result_col60[52] <= result_col60[51];
   result_col60[53] <= result_col60[52];
   result_col60[54] <= result_col60[53];
   result_col60[55] <= result_col60[54];
   result_col60[56] <= result_col60[55];
   result_col60[57] <= result_col60[56];
   result_col60[58] <= result_col60[57];
   result_col60[59] <= result_col60[58];
   result_col60[60] <= result_col60[59];
   result_col60[61] <= result_col60[60];
   result_col60[62] <= result_col60[61];
   result_col60[63] <= result_col60[62];
   result_col60[64] <= result_col60[63];
   result_col60[65] <= result_col60[64];
   result_col60[66] <= result_col60[65];
   result_col60[67] <= result_col60[66];
   result_col60[68] <= result_col60[67];
   result_col60[69] <= result_col60[68];
   result_col60[70] <= result_col60[69];
   result_col60[71] <= result_col60[70];
   result_col60[72] <= result_col60[71];
   result_col60[73] <= result_col60[72];
   result_col60[74] <= result_col60[73];
   result_col60[75] <= result_col60[74];
   result_col60[76] <= result_col60[75];
   result_col60[77] <= result_col60[76];
   result_col60[78] <= result_col60[77];
   result_col60[79] <= result_col60[78];
   result_col60[80] <= result_col60[79];
   result_col60[81] <= result_col60[80];
   result_col60[82] <= result_col60[81];
   result_col60[83] <= result_col60[82];
   result_col60[84] <= result_col60[83];
   result_col60[85] <= result_col60[84];
   result_col60[86] <= result_col60[85];
   result_col60[87] <= result_col60[86];
   result_col60[88] <= result_col60[87];
   result_col60[89] <= result_col60[88];
   result_col60[90] <= result_col60[89];
   result_col60[91] <= result_col60[90];
   result_col60[92] <= result_col60[91];
   result_col60[93] <= result_col60[92];
   result_col60[94] <= result_col60[93];
   result_col60[95] <= result_col60[94];
   result_col60[96] <= result_col60[95];
   result_col60[97] <= result_col60[96];
   result_col60[98] <= result_col60[97];
   result_col60[99] <= result_col60[98];
   result_col60[100] <= result_col60[99];
   result_col60[101] <= result_col60[100];
   result_col60[102] <= result_col60[101];
   result_col60[103] <= result_col60[102];
   result_col60[104] <= result_col60[103];
   result_col60[105] <= result_col60[104];
   result_col60[106] <= result_col60[105];

   result_col61[1] <= data_out_4_61;
   result_col61[2] <= result_col61[1];
   result_col61[3] <= result_col61[2];
   result_col61[4] <= result_col61[3];
   result_col61[5] <= result_col61[4];
   result_col61[6] <= result_col61[5];
   result_col61[7] <= result_col61[6];
   result_col61[8] <= result_col61[7];
   result_col61[9] <= result_col61[8];
   result_col61[10] <= result_col61[9];
   result_col61[11] <= result_col61[10];
   result_col61[12] <= result_col61[11];
   result_col61[13] <= result_col61[12];
   result_col61[14] <= result_col61[13];
   result_col61[15] <= result_col61[14];
   result_col61[16] <= result_col61[15];
   result_col61[17] <= result_col61[16];
   result_col61[18] <= result_col61[17];
   result_col61[19] <= result_col61[18];
   result_col61[20] <= result_col61[19];
   result_col61[21] <= result_col61[20];
   result_col61[22] <= result_col61[21];
   result_col61[23] <= result_col61[22];
   result_col61[24] <= result_col61[23];
   result_col61[25] <= result_col61[24];
   result_col61[26] <= result_col61[25];
   result_col61[27] <= result_col61[26];
   result_col61[28] <= result_col61[27];
   result_col61[29] <= result_col61[28];
   result_col61[30] <= result_col61[29];
   result_col61[31] <= result_col61[30];
   result_col61[32] <= result_col61[31];
   result_col61[33] <= result_col61[32];
   result_col61[34] <= result_col61[33];
   result_col61[35] <= result_col61[34];
   result_col61[36] <= result_col61[35];
   result_col61[37] <= result_col61[36];
   result_col61[38] <= result_col61[37];
   result_col61[39] <= result_col61[38];
   result_col61[40] <= result_col61[39];
   result_col61[41] <= result_col61[40];
   result_col61[42] <= result_col61[41];
   result_col61[43] <= result_col61[42];
   result_col61[44] <= result_col61[43];
   result_col61[45] <= result_col61[44];
   result_col61[46] <= result_col61[45];
   result_col61[47] <= result_col61[46];
   result_col61[48] <= result_col61[47];
   result_col61[49] <= result_col61[48];
   result_col61[50] <= result_col61[49];
   result_col61[51] <= result_col61[50];
   result_col61[52] <= result_col61[51];
   result_col61[53] <= result_col61[52];
   result_col61[54] <= result_col61[53];
   result_col61[55] <= result_col61[54];
   result_col61[56] <= result_col61[55];
   result_col61[57] <= result_col61[56];
   result_col61[58] <= result_col61[57];
   result_col61[59] <= result_col61[58];
   result_col61[60] <= result_col61[59];
   result_col61[61] <= result_col61[60];
   result_col61[62] <= result_col61[61];
   result_col61[63] <= result_col61[62];
   result_col61[64] <= result_col61[63];
   result_col61[65] <= result_col61[64];
   result_col61[66] <= result_col61[65];
   result_col61[67] <= result_col61[66];
   result_col61[68] <= result_col61[67];
   result_col61[69] <= result_col61[68];
   result_col61[70] <= result_col61[69];
   result_col61[71] <= result_col61[70];
   result_col61[72] <= result_col61[71];
   result_col61[73] <= result_col61[72];
   result_col61[74] <= result_col61[73];
   result_col61[75] <= result_col61[74];
   result_col61[76] <= result_col61[75];
   result_col61[77] <= result_col61[76];
   result_col61[78] <= result_col61[77];
   result_col61[79] <= result_col61[78];
   result_col61[80] <= result_col61[79];
   result_col61[81] <= result_col61[80];
   result_col61[82] <= result_col61[81];
   result_col61[83] <= result_col61[82];
   result_col61[84] <= result_col61[83];
   result_col61[85] <= result_col61[84];
   result_col61[86] <= result_col61[85];
   result_col61[87] <= result_col61[86];
   result_col61[88] <= result_col61[87];
   result_col61[89] <= result_col61[88];
   result_col61[90] <= result_col61[89];
   result_col61[91] <= result_col61[90];
   result_col61[92] <= result_col61[91];
   result_col61[93] <= result_col61[92];
   result_col61[94] <= result_col61[93];
   result_col61[95] <= result_col61[94];
   result_col61[96] <= result_col61[95];
   result_col61[97] <= result_col61[96];
   result_col61[98] <= result_col61[97];
   result_col61[99] <= result_col61[98];
   result_col61[100] <= result_col61[99];
   result_col61[101] <= result_col61[100];
   result_col61[102] <= result_col61[101];
   result_col61[103] <= result_col61[102];
   result_col61[104] <= result_col61[103];
   result_col61[105] <= result_col61[104];

   result_col62[1] <= data_out_4_62;
   result_col62[2] <= result_col62[1];
   result_col62[3] <= result_col62[2];
   result_col62[4] <= result_col62[3];
   result_col62[5] <= result_col62[4];
   result_col62[6] <= result_col62[5];
   result_col62[7] <= result_col62[6];
   result_col62[8] <= result_col62[7];
   result_col62[9] <= result_col62[8];
   result_col62[10] <= result_col62[9];
   result_col62[11] <= result_col62[10];
   result_col62[12] <= result_col62[11];
   result_col62[13] <= result_col62[12];
   result_col62[14] <= result_col62[13];
   result_col62[15] <= result_col62[14];
   result_col62[16] <= result_col62[15];
   result_col62[17] <= result_col62[16];
   result_col62[18] <= result_col62[17];
   result_col62[19] <= result_col62[18];
   result_col62[20] <= result_col62[19];
   result_col62[21] <= result_col62[20];
   result_col62[22] <= result_col62[21];
   result_col62[23] <= result_col62[22];
   result_col62[24] <= result_col62[23];
   result_col62[25] <= result_col62[24];
   result_col62[26] <= result_col62[25];
   result_col62[27] <= result_col62[26];
   result_col62[28] <= result_col62[27];
   result_col62[29] <= result_col62[28];
   result_col62[30] <= result_col62[29];
   result_col62[31] <= result_col62[30];
   result_col62[32] <= result_col62[31];
   result_col62[33] <= result_col62[32];
   result_col62[34] <= result_col62[33];
   result_col62[35] <= result_col62[34];
   result_col62[36] <= result_col62[35];
   result_col62[37] <= result_col62[36];
   result_col62[38] <= result_col62[37];
   result_col62[39] <= result_col62[38];
   result_col62[40] <= result_col62[39];
   result_col62[41] <= result_col62[40];
   result_col62[42] <= result_col62[41];
   result_col62[43] <= result_col62[42];
   result_col62[44] <= result_col62[43];
   result_col62[45] <= result_col62[44];
   result_col62[46] <= result_col62[45];
   result_col62[47] <= result_col62[46];
   result_col62[48] <= result_col62[47];
   result_col62[49] <= result_col62[48];
   result_col62[50] <= result_col62[49];
   result_col62[51] <= result_col62[50];
   result_col62[52] <= result_col62[51];
   result_col62[53] <= result_col62[52];
   result_col62[54] <= result_col62[53];
   result_col62[55] <= result_col62[54];
   result_col62[56] <= result_col62[55];
   result_col62[57] <= result_col62[56];
   result_col62[58] <= result_col62[57];
   result_col62[59] <= result_col62[58];
   result_col62[60] <= result_col62[59];
   result_col62[61] <= result_col62[60];
   result_col62[62] <= result_col62[61];
   result_col62[63] <= result_col62[62];
   result_col62[64] <= result_col62[63];
   result_col62[65] <= result_col62[64];
   result_col62[66] <= result_col62[65];
   result_col62[67] <= result_col62[66];
   result_col62[68] <= result_col62[67];
   result_col62[69] <= result_col62[68];
   result_col62[70] <= result_col62[69];
   result_col62[71] <= result_col62[70];
   result_col62[72] <= result_col62[71];
   result_col62[73] <= result_col62[72];
   result_col62[74] <= result_col62[73];
   result_col62[75] <= result_col62[74];
   result_col62[76] <= result_col62[75];
   result_col62[77] <= result_col62[76];
   result_col62[78] <= result_col62[77];
   result_col62[79] <= result_col62[78];
   result_col62[80] <= result_col62[79];
   result_col62[81] <= result_col62[80];
   result_col62[82] <= result_col62[81];
   result_col62[83] <= result_col62[82];
   result_col62[84] <= result_col62[83];
   result_col62[85] <= result_col62[84];
   result_col62[86] <= result_col62[85];
   result_col62[87] <= result_col62[86];
   result_col62[88] <= result_col62[87];
   result_col62[89] <= result_col62[88];
   result_col62[90] <= result_col62[89];
   result_col62[91] <= result_col62[90];
   result_col62[92] <= result_col62[91];
   result_col62[93] <= result_col62[92];
   result_col62[94] <= result_col62[93];
   result_col62[95] <= result_col62[94];
   result_col62[96] <= result_col62[95];
   result_col62[97] <= result_col62[96];
   result_col62[98] <= result_col62[97];
   result_col62[99] <= result_col62[98];
   result_col62[100] <= result_col62[99];
   result_col62[101] <= result_col62[100];
   result_col62[102] <= result_col62[101];
   result_col62[103] <= result_col62[102];
   result_col62[104] <= result_col62[103];

   result_col63[1] <= data_out_4_63;
   result_col63[2] <= result_col63[1];
   result_col63[3] <= result_col63[2];
   result_col63[4] <= result_col63[3];
   result_col63[5] <= result_col63[4];
   result_col63[6] <= result_col63[5];
   result_col63[7] <= result_col63[6];
   result_col63[8] <= result_col63[7];
   result_col63[9] <= result_col63[8];
   result_col63[10] <= result_col63[9];
   result_col63[11] <= result_col63[10];
   result_col63[12] <= result_col63[11];
   result_col63[13] <= result_col63[12];
   result_col63[14] <= result_col63[13];
   result_col63[15] <= result_col63[14];
   result_col63[16] <= result_col63[15];
   result_col63[17] <= result_col63[16];
   result_col63[18] <= result_col63[17];
   result_col63[19] <= result_col63[18];
   result_col63[20] <= result_col63[19];
   result_col63[21] <= result_col63[20];
   result_col63[22] <= result_col63[21];
   result_col63[23] <= result_col63[22];
   result_col63[24] <= result_col63[23];
   result_col63[25] <= result_col63[24];
   result_col63[26] <= result_col63[25];
   result_col63[27] <= result_col63[26];
   result_col63[28] <= result_col63[27];
   result_col63[29] <= result_col63[28];
   result_col63[30] <= result_col63[29];
   result_col63[31] <= result_col63[30];
   result_col63[32] <= result_col63[31];
   result_col63[33] <= result_col63[32];
   result_col63[34] <= result_col63[33];
   result_col63[35] <= result_col63[34];
   result_col63[36] <= result_col63[35];
   result_col63[37] <= result_col63[36];
   result_col63[38] <= result_col63[37];
   result_col63[39] <= result_col63[38];
   result_col63[40] <= result_col63[39];
   result_col63[41] <= result_col63[40];
   result_col63[42] <= result_col63[41];
   result_col63[43] <= result_col63[42];
   result_col63[44] <= result_col63[43];
   result_col63[45] <= result_col63[44];
   result_col63[46] <= result_col63[45];
   result_col63[47] <= result_col63[46];
   result_col63[48] <= result_col63[47];
   result_col63[49] <= result_col63[48];
   result_col63[50] <= result_col63[49];
   result_col63[51] <= result_col63[50];
   result_col63[52] <= result_col63[51];
   result_col63[53] <= result_col63[52];
   result_col63[54] <= result_col63[53];
   result_col63[55] <= result_col63[54];
   result_col63[56] <= result_col63[55];
   result_col63[57] <= result_col63[56];
   result_col63[58] <= result_col63[57];
   result_col63[59] <= result_col63[58];
   result_col63[60] <= result_col63[59];
   result_col63[61] <= result_col63[60];
   result_col63[62] <= result_col63[61];
   result_col63[63] <= result_col63[62];
   result_col63[64] <= result_col63[63];
   result_col63[65] <= result_col63[64];
   result_col63[66] <= result_col63[65];
   result_col63[67] <= result_col63[66];
   result_col63[68] <= result_col63[67];
   result_col63[69] <= result_col63[68];
   result_col63[70] <= result_col63[69];
   result_col63[71] <= result_col63[70];
   result_col63[72] <= result_col63[71];
   result_col63[73] <= result_col63[72];
   result_col63[74] <= result_col63[73];
   result_col63[75] <= result_col63[74];
   result_col63[76] <= result_col63[75];
   result_col63[77] <= result_col63[76];
   result_col63[78] <= result_col63[77];
   result_col63[79] <= result_col63[78];
   result_col63[80] <= result_col63[79];
   result_col63[81] <= result_col63[80];
   result_col63[82] <= result_col63[81];
   result_col63[83] <= result_col63[82];
   result_col63[84] <= result_col63[83];
   result_col63[85] <= result_col63[84];
   result_col63[86] <= result_col63[85];
   result_col63[87] <= result_col63[86];
   result_col63[88] <= result_col63[87];
   result_col63[89] <= result_col63[88];
   result_col63[90] <= result_col63[89];
   result_col63[91] <= result_col63[90];
   result_col63[92] <= result_col63[91];
   result_col63[93] <= result_col63[92];
   result_col63[94] <= result_col63[93];
   result_col63[95] <= result_col63[94];
   result_col63[96] <= result_col63[95];
   result_col63[97] <= result_col63[96];
   result_col63[98] <= result_col63[97];
   result_col63[99] <= result_col63[98];
   result_col63[100] <= result_col63[99];
   result_col63[101] <= result_col63[100];
   result_col63[102] <= result_col63[101];
   result_col63[103] <= result_col63[102];

   result_col64[1] <= data_out_4_64;
   result_col64[2] <= result_col64[1];
   result_col64[3] <= result_col64[2];
   result_col64[4] <= result_col64[3];
   result_col64[5] <= result_col64[4];
   result_col64[6] <= result_col64[5];
   result_col64[7] <= result_col64[6];
   result_col64[8] <= result_col64[7];
   result_col64[9] <= result_col64[8];
   result_col64[10] <= result_col64[9];
   result_col64[11] <= result_col64[10];
   result_col64[12] <= result_col64[11];
   result_col64[13] <= result_col64[12];
   result_col64[14] <= result_col64[13];
   result_col64[15] <= result_col64[14];
   result_col64[16] <= result_col64[15];
   result_col64[17] <= result_col64[16];
   result_col64[18] <= result_col64[17];
   result_col64[19] <= result_col64[18];
   result_col64[20] <= result_col64[19];
   result_col64[21] <= result_col64[20];
   result_col64[22] <= result_col64[21];
   result_col64[23] <= result_col64[22];
   result_col64[24] <= result_col64[23];
   result_col64[25] <= result_col64[24];
   result_col64[26] <= result_col64[25];
   result_col64[27] <= result_col64[26];
   result_col64[28] <= result_col64[27];
   result_col64[29] <= result_col64[28];
   result_col64[30] <= result_col64[29];
   result_col64[31] <= result_col64[30];
   result_col64[32] <= result_col64[31];
   result_col64[33] <= result_col64[32];
   result_col64[34] <= result_col64[33];
   result_col64[35] <= result_col64[34];
   result_col64[36] <= result_col64[35];
   result_col64[37] <= result_col64[36];
   result_col64[38] <= result_col64[37];
   result_col64[39] <= result_col64[38];
   result_col64[40] <= result_col64[39];
   result_col64[41] <= result_col64[40];
   result_col64[42] <= result_col64[41];
   result_col64[43] <= result_col64[42];
   result_col64[44] <= result_col64[43];
   result_col64[45] <= result_col64[44];
   result_col64[46] <= result_col64[45];
   result_col64[47] <= result_col64[46];
   result_col64[48] <= result_col64[47];
   result_col64[49] <= result_col64[48];
   result_col64[50] <= result_col64[49];
   result_col64[51] <= result_col64[50];
   result_col64[52] <= result_col64[51];
   result_col64[53] <= result_col64[52];
   result_col64[54] <= result_col64[53];
   result_col64[55] <= result_col64[54];
   result_col64[56] <= result_col64[55];
   result_col64[57] <= result_col64[56];
   result_col64[58] <= result_col64[57];
   result_col64[59] <= result_col64[58];
   result_col64[60] <= result_col64[59];
   result_col64[61] <= result_col64[60];
   result_col64[62] <= result_col64[61];
   result_col64[63] <= result_col64[62];
   result_col64[64] <= result_col64[63];
   result_col64[65] <= result_col64[64];
   result_col64[66] <= result_col64[65];
   result_col64[67] <= result_col64[66];
   result_col64[68] <= result_col64[67];
   result_col64[69] <= result_col64[68];
   result_col64[70] <= result_col64[69];
   result_col64[71] <= result_col64[70];
   result_col64[72] <= result_col64[71];
   result_col64[73] <= result_col64[72];
   result_col64[74] <= result_col64[73];
   result_col64[75] <= result_col64[74];
   result_col64[76] <= result_col64[75];
   result_col64[77] <= result_col64[76];
   result_col64[78] <= result_col64[77];
   result_col64[79] <= result_col64[78];
   result_col64[80] <= result_col64[79];
   result_col64[81] <= result_col64[80];
   result_col64[82] <= result_col64[81];
   result_col64[83] <= result_col64[82];
   result_col64[84] <= result_col64[83];
   result_col64[85] <= result_col64[84];
   result_col64[86] <= result_col64[85];
   result_col64[87] <= result_col64[86];
   result_col64[88] <= result_col64[87];
   result_col64[89] <= result_col64[88];
   result_col64[90] <= result_col64[89];
   result_col64[91] <= result_col64[90];
   result_col64[92] <= result_col64[91];
   result_col64[93] <= result_col64[92];
   result_col64[94] <= result_col64[93];
   result_col64[95] <= result_col64[94];
   result_col64[96] <= result_col64[95];
   result_col64[97] <= result_col64[96];
   result_col64[98] <= result_col64[97];
   result_col64[99] <= result_col64[98];
   result_col64[100] <= result_col64[99];
   result_col64[101] <= result_col64[100];
   result_col64[102] <= result_col64[101];

   result_col65[1] <= data_out_4_65;
   result_col65[2] <= result_col65[1];
   result_col65[3] <= result_col65[2];
   result_col65[4] <= result_col65[3];
   result_col65[5] <= result_col65[4];
   result_col65[6] <= result_col65[5];
   result_col65[7] <= result_col65[6];
   result_col65[8] <= result_col65[7];
   result_col65[9] <= result_col65[8];
   result_col65[10] <= result_col65[9];
   result_col65[11] <= result_col65[10];
   result_col65[12] <= result_col65[11];
   result_col65[13] <= result_col65[12];
   result_col65[14] <= result_col65[13];
   result_col65[15] <= result_col65[14];
   result_col65[16] <= result_col65[15];
   result_col65[17] <= result_col65[16];
   result_col65[18] <= result_col65[17];
   result_col65[19] <= result_col65[18];
   result_col65[20] <= result_col65[19];
   result_col65[21] <= result_col65[20];
   result_col65[22] <= result_col65[21];
   result_col65[23] <= result_col65[22];
   result_col65[24] <= result_col65[23];
   result_col65[25] <= result_col65[24];
   result_col65[26] <= result_col65[25];
   result_col65[27] <= result_col65[26];
   result_col65[28] <= result_col65[27];
   result_col65[29] <= result_col65[28];
   result_col65[30] <= result_col65[29];
   result_col65[31] <= result_col65[30];
   result_col65[32] <= result_col65[31];
   result_col65[33] <= result_col65[32];
   result_col65[34] <= result_col65[33];
   result_col65[35] <= result_col65[34];
   result_col65[36] <= result_col65[35];
   result_col65[37] <= result_col65[36];
   result_col65[38] <= result_col65[37];
   result_col65[39] <= result_col65[38];
   result_col65[40] <= result_col65[39];
   result_col65[41] <= result_col65[40];
   result_col65[42] <= result_col65[41];
   result_col65[43] <= result_col65[42];
   result_col65[44] <= result_col65[43];
   result_col65[45] <= result_col65[44];
   result_col65[46] <= result_col65[45];
   result_col65[47] <= result_col65[46];
   result_col65[48] <= result_col65[47];
   result_col65[49] <= result_col65[48];
   result_col65[50] <= result_col65[49];
   result_col65[51] <= result_col65[50];
   result_col65[52] <= result_col65[51];
   result_col65[53] <= result_col65[52];
   result_col65[54] <= result_col65[53];
   result_col65[55] <= result_col65[54];
   result_col65[56] <= result_col65[55];
   result_col65[57] <= result_col65[56];
   result_col65[58] <= result_col65[57];
   result_col65[59] <= result_col65[58];
   result_col65[60] <= result_col65[59];
   result_col65[61] <= result_col65[60];
   result_col65[62] <= result_col65[61];
   result_col65[63] <= result_col65[62];
   result_col65[64] <= result_col65[63];
   result_col65[65] <= result_col65[64];
   result_col65[66] <= result_col65[65];
   result_col65[67] <= result_col65[66];
   result_col65[68] <= result_col65[67];
   result_col65[69] <= result_col65[68];
   result_col65[70] <= result_col65[69];
   result_col65[71] <= result_col65[70];
   result_col65[72] <= result_col65[71];
   result_col65[73] <= result_col65[72];
   result_col65[74] <= result_col65[73];
   result_col65[75] <= result_col65[74];
   result_col65[76] <= result_col65[75];
   result_col65[77] <= result_col65[76];
   result_col65[78] <= result_col65[77];
   result_col65[79] <= result_col65[78];
   result_col65[80] <= result_col65[79];
   result_col65[81] <= result_col65[80];
   result_col65[82] <= result_col65[81];
   result_col65[83] <= result_col65[82];
   result_col65[84] <= result_col65[83];
   result_col65[85] <= result_col65[84];
   result_col65[86] <= result_col65[85];
   result_col65[87] <= result_col65[86];
   result_col65[88] <= result_col65[87];
   result_col65[89] <= result_col65[88];
   result_col65[90] <= result_col65[89];
   result_col65[91] <= result_col65[90];
   result_col65[92] <= result_col65[91];
   result_col65[93] <= result_col65[92];
   result_col65[94] <= result_col65[93];
   result_col65[95] <= result_col65[94];
   result_col65[96] <= result_col65[95];
   result_col65[97] <= result_col65[96];
   result_col65[98] <= result_col65[97];
   result_col65[99] <= result_col65[98];
   result_col65[100] <= result_col65[99];
   result_col65[101] <= result_col65[100];

   result_col66[1] <= data_out_4_66;
   result_col66[2] <= result_col66[1];
   result_col66[3] <= result_col66[2];
   result_col66[4] <= result_col66[3];
   result_col66[5] <= result_col66[4];
   result_col66[6] <= result_col66[5];
   result_col66[7] <= result_col66[6];
   result_col66[8] <= result_col66[7];
   result_col66[9] <= result_col66[8];
   result_col66[10] <= result_col66[9];
   result_col66[11] <= result_col66[10];
   result_col66[12] <= result_col66[11];
   result_col66[13] <= result_col66[12];
   result_col66[14] <= result_col66[13];
   result_col66[15] <= result_col66[14];
   result_col66[16] <= result_col66[15];
   result_col66[17] <= result_col66[16];
   result_col66[18] <= result_col66[17];
   result_col66[19] <= result_col66[18];
   result_col66[20] <= result_col66[19];
   result_col66[21] <= result_col66[20];
   result_col66[22] <= result_col66[21];
   result_col66[23] <= result_col66[22];
   result_col66[24] <= result_col66[23];
   result_col66[25] <= result_col66[24];
   result_col66[26] <= result_col66[25];
   result_col66[27] <= result_col66[26];
   result_col66[28] <= result_col66[27];
   result_col66[29] <= result_col66[28];
   result_col66[30] <= result_col66[29];
   result_col66[31] <= result_col66[30];
   result_col66[32] <= result_col66[31];
   result_col66[33] <= result_col66[32];
   result_col66[34] <= result_col66[33];
   result_col66[35] <= result_col66[34];
   result_col66[36] <= result_col66[35];
   result_col66[37] <= result_col66[36];
   result_col66[38] <= result_col66[37];
   result_col66[39] <= result_col66[38];
   result_col66[40] <= result_col66[39];
   result_col66[41] <= result_col66[40];
   result_col66[42] <= result_col66[41];
   result_col66[43] <= result_col66[42];
   result_col66[44] <= result_col66[43];
   result_col66[45] <= result_col66[44];
   result_col66[46] <= result_col66[45];
   result_col66[47] <= result_col66[46];
   result_col66[48] <= result_col66[47];
   result_col66[49] <= result_col66[48];
   result_col66[50] <= result_col66[49];
   result_col66[51] <= result_col66[50];
   result_col66[52] <= result_col66[51];
   result_col66[53] <= result_col66[52];
   result_col66[54] <= result_col66[53];
   result_col66[55] <= result_col66[54];
   result_col66[56] <= result_col66[55];
   result_col66[57] <= result_col66[56];
   result_col66[58] <= result_col66[57];
   result_col66[59] <= result_col66[58];
   result_col66[60] <= result_col66[59];
   result_col66[61] <= result_col66[60];
   result_col66[62] <= result_col66[61];
   result_col66[63] <= result_col66[62];
   result_col66[64] <= result_col66[63];
   result_col66[65] <= result_col66[64];
   result_col66[66] <= result_col66[65];
   result_col66[67] <= result_col66[66];
   result_col66[68] <= result_col66[67];
   result_col66[69] <= result_col66[68];
   result_col66[70] <= result_col66[69];
   result_col66[71] <= result_col66[70];
   result_col66[72] <= result_col66[71];
   result_col66[73] <= result_col66[72];
   result_col66[74] <= result_col66[73];
   result_col66[75] <= result_col66[74];
   result_col66[76] <= result_col66[75];
   result_col66[77] <= result_col66[76];
   result_col66[78] <= result_col66[77];
   result_col66[79] <= result_col66[78];
   result_col66[80] <= result_col66[79];
   result_col66[81] <= result_col66[80];
   result_col66[82] <= result_col66[81];
   result_col66[83] <= result_col66[82];
   result_col66[84] <= result_col66[83];
   result_col66[85] <= result_col66[84];
   result_col66[86] <= result_col66[85];
   result_col66[87] <= result_col66[86];
   result_col66[88] <= result_col66[87];
   result_col66[89] <= result_col66[88];
   result_col66[90] <= result_col66[89];
   result_col66[91] <= result_col66[90];
   result_col66[92] <= result_col66[91];
   result_col66[93] <= result_col66[92];
   result_col66[94] <= result_col66[93];
   result_col66[95] <= result_col66[94];
   result_col66[96] <= result_col66[95];
   result_col66[97] <= result_col66[96];
   result_col66[98] <= result_col66[97];
   result_col66[99] <= result_col66[98];
   result_col66[100] <= result_col66[99];

   result_col67[1] <= data_out_4_67;
   result_col67[2] <= result_col67[1];
   result_col67[3] <= result_col67[2];
   result_col67[4] <= result_col67[3];
   result_col67[5] <= result_col67[4];
   result_col67[6] <= result_col67[5];
   result_col67[7] <= result_col67[6];
   result_col67[8] <= result_col67[7];
   result_col67[9] <= result_col67[8];
   result_col67[10] <= result_col67[9];
   result_col67[11] <= result_col67[10];
   result_col67[12] <= result_col67[11];
   result_col67[13] <= result_col67[12];
   result_col67[14] <= result_col67[13];
   result_col67[15] <= result_col67[14];
   result_col67[16] <= result_col67[15];
   result_col67[17] <= result_col67[16];
   result_col67[18] <= result_col67[17];
   result_col67[19] <= result_col67[18];
   result_col67[20] <= result_col67[19];
   result_col67[21] <= result_col67[20];
   result_col67[22] <= result_col67[21];
   result_col67[23] <= result_col67[22];
   result_col67[24] <= result_col67[23];
   result_col67[25] <= result_col67[24];
   result_col67[26] <= result_col67[25];
   result_col67[27] <= result_col67[26];
   result_col67[28] <= result_col67[27];
   result_col67[29] <= result_col67[28];
   result_col67[30] <= result_col67[29];
   result_col67[31] <= result_col67[30];
   result_col67[32] <= result_col67[31];
   result_col67[33] <= result_col67[32];
   result_col67[34] <= result_col67[33];
   result_col67[35] <= result_col67[34];
   result_col67[36] <= result_col67[35];
   result_col67[37] <= result_col67[36];
   result_col67[38] <= result_col67[37];
   result_col67[39] <= result_col67[38];
   result_col67[40] <= result_col67[39];
   result_col67[41] <= result_col67[40];
   result_col67[42] <= result_col67[41];
   result_col67[43] <= result_col67[42];
   result_col67[44] <= result_col67[43];
   result_col67[45] <= result_col67[44];
   result_col67[46] <= result_col67[45];
   result_col67[47] <= result_col67[46];
   result_col67[48] <= result_col67[47];
   result_col67[49] <= result_col67[48];
   result_col67[50] <= result_col67[49];
   result_col67[51] <= result_col67[50];
   result_col67[52] <= result_col67[51];
   result_col67[53] <= result_col67[52];
   result_col67[54] <= result_col67[53];
   result_col67[55] <= result_col67[54];
   result_col67[56] <= result_col67[55];
   result_col67[57] <= result_col67[56];
   result_col67[58] <= result_col67[57];
   result_col67[59] <= result_col67[58];
   result_col67[60] <= result_col67[59];
   result_col67[61] <= result_col67[60];
   result_col67[62] <= result_col67[61];
   result_col67[63] <= result_col67[62];
   result_col67[64] <= result_col67[63];
   result_col67[65] <= result_col67[64];
   result_col67[66] <= result_col67[65];
   result_col67[67] <= result_col67[66];
   result_col67[68] <= result_col67[67];
   result_col67[69] <= result_col67[68];
   result_col67[70] <= result_col67[69];
   result_col67[71] <= result_col67[70];
   result_col67[72] <= result_col67[71];
   result_col67[73] <= result_col67[72];
   result_col67[74] <= result_col67[73];
   result_col67[75] <= result_col67[74];
   result_col67[76] <= result_col67[75];
   result_col67[77] <= result_col67[76];
   result_col67[78] <= result_col67[77];
   result_col67[79] <= result_col67[78];
   result_col67[80] <= result_col67[79];
   result_col67[81] <= result_col67[80];
   result_col67[82] <= result_col67[81];
   result_col67[83] <= result_col67[82];
   result_col67[84] <= result_col67[83];
   result_col67[85] <= result_col67[84];
   result_col67[86] <= result_col67[85];
   result_col67[87] <= result_col67[86];
   result_col67[88] <= result_col67[87];
   result_col67[89] <= result_col67[88];
   result_col67[90] <= result_col67[89];
   result_col67[91] <= result_col67[90];
   result_col67[92] <= result_col67[91];
   result_col67[93] <= result_col67[92];
   result_col67[94] <= result_col67[93];
   result_col67[95] <= result_col67[94];
   result_col67[96] <= result_col67[95];
   result_col67[97] <= result_col67[96];
   result_col67[98] <= result_col67[97];
   result_col67[99] <= result_col67[98];

   result_col68[1] <= data_out_4_68;
   result_col68[2] <= result_col68[1];
   result_col68[3] <= result_col68[2];
   result_col68[4] <= result_col68[3];
   result_col68[5] <= result_col68[4];
   result_col68[6] <= result_col68[5];
   result_col68[7] <= result_col68[6];
   result_col68[8] <= result_col68[7];
   result_col68[9] <= result_col68[8];
   result_col68[10] <= result_col68[9];
   result_col68[11] <= result_col68[10];
   result_col68[12] <= result_col68[11];
   result_col68[13] <= result_col68[12];
   result_col68[14] <= result_col68[13];
   result_col68[15] <= result_col68[14];
   result_col68[16] <= result_col68[15];
   result_col68[17] <= result_col68[16];
   result_col68[18] <= result_col68[17];
   result_col68[19] <= result_col68[18];
   result_col68[20] <= result_col68[19];
   result_col68[21] <= result_col68[20];
   result_col68[22] <= result_col68[21];
   result_col68[23] <= result_col68[22];
   result_col68[24] <= result_col68[23];
   result_col68[25] <= result_col68[24];
   result_col68[26] <= result_col68[25];
   result_col68[27] <= result_col68[26];
   result_col68[28] <= result_col68[27];
   result_col68[29] <= result_col68[28];
   result_col68[30] <= result_col68[29];
   result_col68[31] <= result_col68[30];
   result_col68[32] <= result_col68[31];
   result_col68[33] <= result_col68[32];
   result_col68[34] <= result_col68[33];
   result_col68[35] <= result_col68[34];
   result_col68[36] <= result_col68[35];
   result_col68[37] <= result_col68[36];
   result_col68[38] <= result_col68[37];
   result_col68[39] <= result_col68[38];
   result_col68[40] <= result_col68[39];
   result_col68[41] <= result_col68[40];
   result_col68[42] <= result_col68[41];
   result_col68[43] <= result_col68[42];
   result_col68[44] <= result_col68[43];
   result_col68[45] <= result_col68[44];
   result_col68[46] <= result_col68[45];
   result_col68[47] <= result_col68[46];
   result_col68[48] <= result_col68[47];
   result_col68[49] <= result_col68[48];
   result_col68[50] <= result_col68[49];
   result_col68[51] <= result_col68[50];
   result_col68[52] <= result_col68[51];
   result_col68[53] <= result_col68[52];
   result_col68[54] <= result_col68[53];
   result_col68[55] <= result_col68[54];
   result_col68[56] <= result_col68[55];
   result_col68[57] <= result_col68[56];
   result_col68[58] <= result_col68[57];
   result_col68[59] <= result_col68[58];
   result_col68[60] <= result_col68[59];
   result_col68[61] <= result_col68[60];
   result_col68[62] <= result_col68[61];
   result_col68[63] <= result_col68[62];
   result_col68[64] <= result_col68[63];
   result_col68[65] <= result_col68[64];
   result_col68[66] <= result_col68[65];
   result_col68[67] <= result_col68[66];
   result_col68[68] <= result_col68[67];
   result_col68[69] <= result_col68[68];
   result_col68[70] <= result_col68[69];
   result_col68[71] <= result_col68[70];
   result_col68[72] <= result_col68[71];
   result_col68[73] <= result_col68[72];
   result_col68[74] <= result_col68[73];
   result_col68[75] <= result_col68[74];
   result_col68[76] <= result_col68[75];
   result_col68[77] <= result_col68[76];
   result_col68[78] <= result_col68[77];
   result_col68[79] <= result_col68[78];
   result_col68[80] <= result_col68[79];
   result_col68[81] <= result_col68[80];
   result_col68[82] <= result_col68[81];
   result_col68[83] <= result_col68[82];
   result_col68[84] <= result_col68[83];
   result_col68[85] <= result_col68[84];
   result_col68[86] <= result_col68[85];
   result_col68[87] <= result_col68[86];
   result_col68[88] <= result_col68[87];
   result_col68[89] <= result_col68[88];
   result_col68[90] <= result_col68[89];
   result_col68[91] <= result_col68[90];
   result_col68[92] <= result_col68[91];
   result_col68[93] <= result_col68[92];
   result_col68[94] <= result_col68[93];
   result_col68[95] <= result_col68[94];
   result_col68[96] <= result_col68[95];
   result_col68[97] <= result_col68[96];
   result_col68[98] <= result_col68[97];

   result_col69[1] <= data_out_4_69;
   result_col69[2] <= result_col69[1];
   result_col69[3] <= result_col69[2];
   result_col69[4] <= result_col69[3];
   result_col69[5] <= result_col69[4];
   result_col69[6] <= result_col69[5];
   result_col69[7] <= result_col69[6];
   result_col69[8] <= result_col69[7];
   result_col69[9] <= result_col69[8];
   result_col69[10] <= result_col69[9];
   result_col69[11] <= result_col69[10];
   result_col69[12] <= result_col69[11];
   result_col69[13] <= result_col69[12];
   result_col69[14] <= result_col69[13];
   result_col69[15] <= result_col69[14];
   result_col69[16] <= result_col69[15];
   result_col69[17] <= result_col69[16];
   result_col69[18] <= result_col69[17];
   result_col69[19] <= result_col69[18];
   result_col69[20] <= result_col69[19];
   result_col69[21] <= result_col69[20];
   result_col69[22] <= result_col69[21];
   result_col69[23] <= result_col69[22];
   result_col69[24] <= result_col69[23];
   result_col69[25] <= result_col69[24];
   result_col69[26] <= result_col69[25];
   result_col69[27] <= result_col69[26];
   result_col69[28] <= result_col69[27];
   result_col69[29] <= result_col69[28];
   result_col69[30] <= result_col69[29];
   result_col69[31] <= result_col69[30];
   result_col69[32] <= result_col69[31];
   result_col69[33] <= result_col69[32];
   result_col69[34] <= result_col69[33];
   result_col69[35] <= result_col69[34];
   result_col69[36] <= result_col69[35];
   result_col69[37] <= result_col69[36];
   result_col69[38] <= result_col69[37];
   result_col69[39] <= result_col69[38];
   result_col69[40] <= result_col69[39];
   result_col69[41] <= result_col69[40];
   result_col69[42] <= result_col69[41];
   result_col69[43] <= result_col69[42];
   result_col69[44] <= result_col69[43];
   result_col69[45] <= result_col69[44];
   result_col69[46] <= result_col69[45];
   result_col69[47] <= result_col69[46];
   result_col69[48] <= result_col69[47];
   result_col69[49] <= result_col69[48];
   result_col69[50] <= result_col69[49];
   result_col69[51] <= result_col69[50];
   result_col69[52] <= result_col69[51];
   result_col69[53] <= result_col69[52];
   result_col69[54] <= result_col69[53];
   result_col69[55] <= result_col69[54];
   result_col69[56] <= result_col69[55];
   result_col69[57] <= result_col69[56];
   result_col69[58] <= result_col69[57];
   result_col69[59] <= result_col69[58];
   result_col69[60] <= result_col69[59];
   result_col69[61] <= result_col69[60];
   result_col69[62] <= result_col69[61];
   result_col69[63] <= result_col69[62];
   result_col69[64] <= result_col69[63];
   result_col69[65] <= result_col69[64];
   result_col69[66] <= result_col69[65];
   result_col69[67] <= result_col69[66];
   result_col69[68] <= result_col69[67];
   result_col69[69] <= result_col69[68];
   result_col69[70] <= result_col69[69];
   result_col69[71] <= result_col69[70];
   result_col69[72] <= result_col69[71];
   result_col69[73] <= result_col69[72];
   result_col69[74] <= result_col69[73];
   result_col69[75] <= result_col69[74];
   result_col69[76] <= result_col69[75];
   result_col69[77] <= result_col69[76];
   result_col69[78] <= result_col69[77];
   result_col69[79] <= result_col69[78];
   result_col69[80] <= result_col69[79];
   result_col69[81] <= result_col69[80];
   result_col69[82] <= result_col69[81];
   result_col69[83] <= result_col69[82];
   result_col69[84] <= result_col69[83];
   result_col69[85] <= result_col69[84];
   result_col69[86] <= result_col69[85];
   result_col69[87] <= result_col69[86];
   result_col69[88] <= result_col69[87];
   result_col69[89] <= result_col69[88];
   result_col69[90] <= result_col69[89];
   result_col69[91] <= result_col69[90];
   result_col69[92] <= result_col69[91];
   result_col69[93] <= result_col69[92];
   result_col69[94] <= result_col69[93];
   result_col69[95] <= result_col69[94];
   result_col69[96] <= result_col69[95];
   result_col69[97] <= result_col69[96];

   result_col70[1] <= data_out_4_70;
   result_col70[2] <= result_col70[1];
   result_col70[3] <= result_col70[2];
   result_col70[4] <= result_col70[3];
   result_col70[5] <= result_col70[4];
   result_col70[6] <= result_col70[5];
   result_col70[7] <= result_col70[6];
   result_col70[8] <= result_col70[7];
   result_col70[9] <= result_col70[8];
   result_col70[10] <= result_col70[9];
   result_col70[11] <= result_col70[10];
   result_col70[12] <= result_col70[11];
   result_col70[13] <= result_col70[12];
   result_col70[14] <= result_col70[13];
   result_col70[15] <= result_col70[14];
   result_col70[16] <= result_col70[15];
   result_col70[17] <= result_col70[16];
   result_col70[18] <= result_col70[17];
   result_col70[19] <= result_col70[18];
   result_col70[20] <= result_col70[19];
   result_col70[21] <= result_col70[20];
   result_col70[22] <= result_col70[21];
   result_col70[23] <= result_col70[22];
   result_col70[24] <= result_col70[23];
   result_col70[25] <= result_col70[24];
   result_col70[26] <= result_col70[25];
   result_col70[27] <= result_col70[26];
   result_col70[28] <= result_col70[27];
   result_col70[29] <= result_col70[28];
   result_col70[30] <= result_col70[29];
   result_col70[31] <= result_col70[30];
   result_col70[32] <= result_col70[31];
   result_col70[33] <= result_col70[32];
   result_col70[34] <= result_col70[33];
   result_col70[35] <= result_col70[34];
   result_col70[36] <= result_col70[35];
   result_col70[37] <= result_col70[36];
   result_col70[38] <= result_col70[37];
   result_col70[39] <= result_col70[38];
   result_col70[40] <= result_col70[39];
   result_col70[41] <= result_col70[40];
   result_col70[42] <= result_col70[41];
   result_col70[43] <= result_col70[42];
   result_col70[44] <= result_col70[43];
   result_col70[45] <= result_col70[44];
   result_col70[46] <= result_col70[45];
   result_col70[47] <= result_col70[46];
   result_col70[48] <= result_col70[47];
   result_col70[49] <= result_col70[48];
   result_col70[50] <= result_col70[49];
   result_col70[51] <= result_col70[50];
   result_col70[52] <= result_col70[51];
   result_col70[53] <= result_col70[52];
   result_col70[54] <= result_col70[53];
   result_col70[55] <= result_col70[54];
   result_col70[56] <= result_col70[55];
   result_col70[57] <= result_col70[56];
   result_col70[58] <= result_col70[57];
   result_col70[59] <= result_col70[58];
   result_col70[60] <= result_col70[59];
   result_col70[61] <= result_col70[60];
   result_col70[62] <= result_col70[61];
   result_col70[63] <= result_col70[62];
   result_col70[64] <= result_col70[63];
   result_col70[65] <= result_col70[64];
   result_col70[66] <= result_col70[65];
   result_col70[67] <= result_col70[66];
   result_col70[68] <= result_col70[67];
   result_col70[69] <= result_col70[68];
   result_col70[70] <= result_col70[69];
   result_col70[71] <= result_col70[70];
   result_col70[72] <= result_col70[71];
   result_col70[73] <= result_col70[72];
   result_col70[74] <= result_col70[73];
   result_col70[75] <= result_col70[74];
   result_col70[76] <= result_col70[75];
   result_col70[77] <= result_col70[76];
   result_col70[78] <= result_col70[77];
   result_col70[79] <= result_col70[78];
   result_col70[80] <= result_col70[79];
   result_col70[81] <= result_col70[80];
   result_col70[82] <= result_col70[81];
   result_col70[83] <= result_col70[82];
   result_col70[84] <= result_col70[83];
   result_col70[85] <= result_col70[84];
   result_col70[86] <= result_col70[85];
   result_col70[87] <= result_col70[86];
   result_col70[88] <= result_col70[87];
   result_col70[89] <= result_col70[88];
   result_col70[90] <= result_col70[89];
   result_col70[91] <= result_col70[90];
   result_col70[92] <= result_col70[91];
   result_col70[93] <= result_col70[92];
   result_col70[94] <= result_col70[93];
   result_col70[95] <= result_col70[94];
   result_col70[96] <= result_col70[95];

   result_col71[1] <= data_out_4_71;
   result_col71[2] <= result_col71[1];
   result_col71[3] <= result_col71[2];
   result_col71[4] <= result_col71[3];
   result_col71[5] <= result_col71[4];
   result_col71[6] <= result_col71[5];
   result_col71[7] <= result_col71[6];
   result_col71[8] <= result_col71[7];
   result_col71[9] <= result_col71[8];
   result_col71[10] <= result_col71[9];
   result_col71[11] <= result_col71[10];
   result_col71[12] <= result_col71[11];
   result_col71[13] <= result_col71[12];
   result_col71[14] <= result_col71[13];
   result_col71[15] <= result_col71[14];
   result_col71[16] <= result_col71[15];
   result_col71[17] <= result_col71[16];
   result_col71[18] <= result_col71[17];
   result_col71[19] <= result_col71[18];
   result_col71[20] <= result_col71[19];
   result_col71[21] <= result_col71[20];
   result_col71[22] <= result_col71[21];
   result_col71[23] <= result_col71[22];
   result_col71[24] <= result_col71[23];
   result_col71[25] <= result_col71[24];
   result_col71[26] <= result_col71[25];
   result_col71[27] <= result_col71[26];
   result_col71[28] <= result_col71[27];
   result_col71[29] <= result_col71[28];
   result_col71[30] <= result_col71[29];
   result_col71[31] <= result_col71[30];
   result_col71[32] <= result_col71[31];
   result_col71[33] <= result_col71[32];
   result_col71[34] <= result_col71[33];
   result_col71[35] <= result_col71[34];
   result_col71[36] <= result_col71[35];
   result_col71[37] <= result_col71[36];
   result_col71[38] <= result_col71[37];
   result_col71[39] <= result_col71[38];
   result_col71[40] <= result_col71[39];
   result_col71[41] <= result_col71[40];
   result_col71[42] <= result_col71[41];
   result_col71[43] <= result_col71[42];
   result_col71[44] <= result_col71[43];
   result_col71[45] <= result_col71[44];
   result_col71[46] <= result_col71[45];
   result_col71[47] <= result_col71[46];
   result_col71[48] <= result_col71[47];
   result_col71[49] <= result_col71[48];
   result_col71[50] <= result_col71[49];
   result_col71[51] <= result_col71[50];
   result_col71[52] <= result_col71[51];
   result_col71[53] <= result_col71[52];
   result_col71[54] <= result_col71[53];
   result_col71[55] <= result_col71[54];
   result_col71[56] <= result_col71[55];
   result_col71[57] <= result_col71[56];
   result_col71[58] <= result_col71[57];
   result_col71[59] <= result_col71[58];
   result_col71[60] <= result_col71[59];
   result_col71[61] <= result_col71[60];
   result_col71[62] <= result_col71[61];
   result_col71[63] <= result_col71[62];
   result_col71[64] <= result_col71[63];
   result_col71[65] <= result_col71[64];
   result_col71[66] <= result_col71[65];
   result_col71[67] <= result_col71[66];
   result_col71[68] <= result_col71[67];
   result_col71[69] <= result_col71[68];
   result_col71[70] <= result_col71[69];
   result_col71[71] <= result_col71[70];
   result_col71[72] <= result_col71[71];
   result_col71[73] <= result_col71[72];
   result_col71[74] <= result_col71[73];
   result_col71[75] <= result_col71[74];
   result_col71[76] <= result_col71[75];
   result_col71[77] <= result_col71[76];
   result_col71[78] <= result_col71[77];
   result_col71[79] <= result_col71[78];
   result_col71[80] <= result_col71[79];
   result_col71[81] <= result_col71[80];
   result_col71[82] <= result_col71[81];
   result_col71[83] <= result_col71[82];
   result_col71[84] <= result_col71[83];
   result_col71[85] <= result_col71[84];
   result_col71[86] <= result_col71[85];
   result_col71[87] <= result_col71[86];
   result_col71[88] <= result_col71[87];
   result_col71[89] <= result_col71[88];
   result_col71[90] <= result_col71[89];
   result_col71[91] <= result_col71[90];
   result_col71[92] <= result_col71[91];
   result_col71[93] <= result_col71[92];
   result_col71[94] <= result_col71[93];
   result_col71[95] <= result_col71[94];

   result_col72[1] <= data_out_4_72;
   result_col72[2] <= result_col72[1];
   result_col72[3] <= result_col72[2];
   result_col72[4] <= result_col72[3];
   result_col72[5] <= result_col72[4];
   result_col72[6] <= result_col72[5];
   result_col72[7] <= result_col72[6];
   result_col72[8] <= result_col72[7];
   result_col72[9] <= result_col72[8];
   result_col72[10] <= result_col72[9];
   result_col72[11] <= result_col72[10];
   result_col72[12] <= result_col72[11];
   result_col72[13] <= result_col72[12];
   result_col72[14] <= result_col72[13];
   result_col72[15] <= result_col72[14];
   result_col72[16] <= result_col72[15];
   result_col72[17] <= result_col72[16];
   result_col72[18] <= result_col72[17];
   result_col72[19] <= result_col72[18];
   result_col72[20] <= result_col72[19];
   result_col72[21] <= result_col72[20];
   result_col72[22] <= result_col72[21];
   result_col72[23] <= result_col72[22];
   result_col72[24] <= result_col72[23];
   result_col72[25] <= result_col72[24];
   result_col72[26] <= result_col72[25];
   result_col72[27] <= result_col72[26];
   result_col72[28] <= result_col72[27];
   result_col72[29] <= result_col72[28];
   result_col72[30] <= result_col72[29];
   result_col72[31] <= result_col72[30];
   result_col72[32] <= result_col72[31];
   result_col72[33] <= result_col72[32];
   result_col72[34] <= result_col72[33];
   result_col72[35] <= result_col72[34];
   result_col72[36] <= result_col72[35];
   result_col72[37] <= result_col72[36];
   result_col72[38] <= result_col72[37];
   result_col72[39] <= result_col72[38];
   result_col72[40] <= result_col72[39];
   result_col72[41] <= result_col72[40];
   result_col72[42] <= result_col72[41];
   result_col72[43] <= result_col72[42];
   result_col72[44] <= result_col72[43];
   result_col72[45] <= result_col72[44];
   result_col72[46] <= result_col72[45];
   result_col72[47] <= result_col72[46];
   result_col72[48] <= result_col72[47];
   result_col72[49] <= result_col72[48];
   result_col72[50] <= result_col72[49];
   result_col72[51] <= result_col72[50];
   result_col72[52] <= result_col72[51];
   result_col72[53] <= result_col72[52];
   result_col72[54] <= result_col72[53];
   result_col72[55] <= result_col72[54];
   result_col72[56] <= result_col72[55];
   result_col72[57] <= result_col72[56];
   result_col72[58] <= result_col72[57];
   result_col72[59] <= result_col72[58];
   result_col72[60] <= result_col72[59];
   result_col72[61] <= result_col72[60];
   result_col72[62] <= result_col72[61];
   result_col72[63] <= result_col72[62];
   result_col72[64] <= result_col72[63];
   result_col72[65] <= result_col72[64];
   result_col72[66] <= result_col72[65];
   result_col72[67] <= result_col72[66];
   result_col72[68] <= result_col72[67];
   result_col72[69] <= result_col72[68];
   result_col72[70] <= result_col72[69];
   result_col72[71] <= result_col72[70];
   result_col72[72] <= result_col72[71];
   result_col72[73] <= result_col72[72];
   result_col72[74] <= result_col72[73];
   result_col72[75] <= result_col72[74];
   result_col72[76] <= result_col72[75];
   result_col72[77] <= result_col72[76];
   result_col72[78] <= result_col72[77];
   result_col72[79] <= result_col72[78];
   result_col72[80] <= result_col72[79];
   result_col72[81] <= result_col72[80];
   result_col72[82] <= result_col72[81];
   result_col72[83] <= result_col72[82];
   result_col72[84] <= result_col72[83];
   result_col72[85] <= result_col72[84];
   result_col72[86] <= result_col72[85];
   result_col72[87] <= result_col72[86];
   result_col72[88] <= result_col72[87];
   result_col72[89] <= result_col72[88];
   result_col72[90] <= result_col72[89];
   result_col72[91] <= result_col72[90];
   result_col72[92] <= result_col72[91];
   result_col72[93] <= result_col72[92];
   result_col72[94] <= result_col72[93];

   result_col73[1] <= data_out_4_73;
   result_col73[2] <= result_col73[1];
   result_col73[3] <= result_col73[2];
   result_col73[4] <= result_col73[3];
   result_col73[5] <= result_col73[4];
   result_col73[6] <= result_col73[5];
   result_col73[7] <= result_col73[6];
   result_col73[8] <= result_col73[7];
   result_col73[9] <= result_col73[8];
   result_col73[10] <= result_col73[9];
   result_col73[11] <= result_col73[10];
   result_col73[12] <= result_col73[11];
   result_col73[13] <= result_col73[12];
   result_col73[14] <= result_col73[13];
   result_col73[15] <= result_col73[14];
   result_col73[16] <= result_col73[15];
   result_col73[17] <= result_col73[16];
   result_col73[18] <= result_col73[17];
   result_col73[19] <= result_col73[18];
   result_col73[20] <= result_col73[19];
   result_col73[21] <= result_col73[20];
   result_col73[22] <= result_col73[21];
   result_col73[23] <= result_col73[22];
   result_col73[24] <= result_col73[23];
   result_col73[25] <= result_col73[24];
   result_col73[26] <= result_col73[25];
   result_col73[27] <= result_col73[26];
   result_col73[28] <= result_col73[27];
   result_col73[29] <= result_col73[28];
   result_col73[30] <= result_col73[29];
   result_col73[31] <= result_col73[30];
   result_col73[32] <= result_col73[31];
   result_col73[33] <= result_col73[32];
   result_col73[34] <= result_col73[33];
   result_col73[35] <= result_col73[34];
   result_col73[36] <= result_col73[35];
   result_col73[37] <= result_col73[36];
   result_col73[38] <= result_col73[37];
   result_col73[39] <= result_col73[38];
   result_col73[40] <= result_col73[39];
   result_col73[41] <= result_col73[40];
   result_col73[42] <= result_col73[41];
   result_col73[43] <= result_col73[42];
   result_col73[44] <= result_col73[43];
   result_col73[45] <= result_col73[44];
   result_col73[46] <= result_col73[45];
   result_col73[47] <= result_col73[46];
   result_col73[48] <= result_col73[47];
   result_col73[49] <= result_col73[48];
   result_col73[50] <= result_col73[49];
   result_col73[51] <= result_col73[50];
   result_col73[52] <= result_col73[51];
   result_col73[53] <= result_col73[52];
   result_col73[54] <= result_col73[53];
   result_col73[55] <= result_col73[54];
   result_col73[56] <= result_col73[55];
   result_col73[57] <= result_col73[56];
   result_col73[58] <= result_col73[57];
   result_col73[59] <= result_col73[58];
   result_col73[60] <= result_col73[59];
   result_col73[61] <= result_col73[60];
   result_col73[62] <= result_col73[61];
   result_col73[63] <= result_col73[62];
   result_col73[64] <= result_col73[63];
   result_col73[65] <= result_col73[64];
   result_col73[66] <= result_col73[65];
   result_col73[67] <= result_col73[66];
   result_col73[68] <= result_col73[67];
   result_col73[69] <= result_col73[68];
   result_col73[70] <= result_col73[69];
   result_col73[71] <= result_col73[70];
   result_col73[72] <= result_col73[71];
   result_col73[73] <= result_col73[72];
   result_col73[74] <= result_col73[73];
   result_col73[75] <= result_col73[74];
   result_col73[76] <= result_col73[75];
   result_col73[77] <= result_col73[76];
   result_col73[78] <= result_col73[77];
   result_col73[79] <= result_col73[78];
   result_col73[80] <= result_col73[79];
   result_col73[81] <= result_col73[80];
   result_col73[82] <= result_col73[81];
   result_col73[83] <= result_col73[82];
   result_col73[84] <= result_col73[83];
   result_col73[85] <= result_col73[84];
   result_col73[86] <= result_col73[85];
   result_col73[87] <= result_col73[86];
   result_col73[88] <= result_col73[87];
   result_col73[89] <= result_col73[88];
   result_col73[90] <= result_col73[89];
   result_col73[91] <= result_col73[90];
   result_col73[92] <= result_col73[91];
   result_col73[93] <= result_col73[92];

   result_col74[1] <= data_out_4_74;
   result_col74[2] <= result_col74[1];
   result_col74[3] <= result_col74[2];
   result_col74[4] <= result_col74[3];
   result_col74[5] <= result_col74[4];
   result_col74[6] <= result_col74[5];
   result_col74[7] <= result_col74[6];
   result_col74[8] <= result_col74[7];
   result_col74[9] <= result_col74[8];
   result_col74[10] <= result_col74[9];
   result_col74[11] <= result_col74[10];
   result_col74[12] <= result_col74[11];
   result_col74[13] <= result_col74[12];
   result_col74[14] <= result_col74[13];
   result_col74[15] <= result_col74[14];
   result_col74[16] <= result_col74[15];
   result_col74[17] <= result_col74[16];
   result_col74[18] <= result_col74[17];
   result_col74[19] <= result_col74[18];
   result_col74[20] <= result_col74[19];
   result_col74[21] <= result_col74[20];
   result_col74[22] <= result_col74[21];
   result_col74[23] <= result_col74[22];
   result_col74[24] <= result_col74[23];
   result_col74[25] <= result_col74[24];
   result_col74[26] <= result_col74[25];
   result_col74[27] <= result_col74[26];
   result_col74[28] <= result_col74[27];
   result_col74[29] <= result_col74[28];
   result_col74[30] <= result_col74[29];
   result_col74[31] <= result_col74[30];
   result_col74[32] <= result_col74[31];
   result_col74[33] <= result_col74[32];
   result_col74[34] <= result_col74[33];
   result_col74[35] <= result_col74[34];
   result_col74[36] <= result_col74[35];
   result_col74[37] <= result_col74[36];
   result_col74[38] <= result_col74[37];
   result_col74[39] <= result_col74[38];
   result_col74[40] <= result_col74[39];
   result_col74[41] <= result_col74[40];
   result_col74[42] <= result_col74[41];
   result_col74[43] <= result_col74[42];
   result_col74[44] <= result_col74[43];
   result_col74[45] <= result_col74[44];
   result_col74[46] <= result_col74[45];
   result_col74[47] <= result_col74[46];
   result_col74[48] <= result_col74[47];
   result_col74[49] <= result_col74[48];
   result_col74[50] <= result_col74[49];
   result_col74[51] <= result_col74[50];
   result_col74[52] <= result_col74[51];
   result_col74[53] <= result_col74[52];
   result_col74[54] <= result_col74[53];
   result_col74[55] <= result_col74[54];
   result_col74[56] <= result_col74[55];
   result_col74[57] <= result_col74[56];
   result_col74[58] <= result_col74[57];
   result_col74[59] <= result_col74[58];
   result_col74[60] <= result_col74[59];
   result_col74[61] <= result_col74[60];
   result_col74[62] <= result_col74[61];
   result_col74[63] <= result_col74[62];
   result_col74[64] <= result_col74[63];
   result_col74[65] <= result_col74[64];
   result_col74[66] <= result_col74[65];
   result_col74[67] <= result_col74[66];
   result_col74[68] <= result_col74[67];
   result_col74[69] <= result_col74[68];
   result_col74[70] <= result_col74[69];
   result_col74[71] <= result_col74[70];
   result_col74[72] <= result_col74[71];
   result_col74[73] <= result_col74[72];
   result_col74[74] <= result_col74[73];
   result_col74[75] <= result_col74[74];
   result_col74[76] <= result_col74[75];
   result_col74[77] <= result_col74[76];
   result_col74[78] <= result_col74[77];
   result_col74[79] <= result_col74[78];
   result_col74[80] <= result_col74[79];
   result_col74[81] <= result_col74[80];
   result_col74[82] <= result_col74[81];
   result_col74[83] <= result_col74[82];
   result_col74[84] <= result_col74[83];
   result_col74[85] <= result_col74[84];
   result_col74[86] <= result_col74[85];
   result_col74[87] <= result_col74[86];
   result_col74[88] <= result_col74[87];
   result_col74[89] <= result_col74[88];
   result_col74[90] <= result_col74[89];
   result_col74[91] <= result_col74[90];
   result_col74[92] <= result_col74[91];

   result_col75[1] <= data_out_4_75;
   result_col75[2] <= result_col75[1];
   result_col75[3] <= result_col75[2];
   result_col75[4] <= result_col75[3];
   result_col75[5] <= result_col75[4];
   result_col75[6] <= result_col75[5];
   result_col75[7] <= result_col75[6];
   result_col75[8] <= result_col75[7];
   result_col75[9] <= result_col75[8];
   result_col75[10] <= result_col75[9];
   result_col75[11] <= result_col75[10];
   result_col75[12] <= result_col75[11];
   result_col75[13] <= result_col75[12];
   result_col75[14] <= result_col75[13];
   result_col75[15] <= result_col75[14];
   result_col75[16] <= result_col75[15];
   result_col75[17] <= result_col75[16];
   result_col75[18] <= result_col75[17];
   result_col75[19] <= result_col75[18];
   result_col75[20] <= result_col75[19];
   result_col75[21] <= result_col75[20];
   result_col75[22] <= result_col75[21];
   result_col75[23] <= result_col75[22];
   result_col75[24] <= result_col75[23];
   result_col75[25] <= result_col75[24];
   result_col75[26] <= result_col75[25];
   result_col75[27] <= result_col75[26];
   result_col75[28] <= result_col75[27];
   result_col75[29] <= result_col75[28];
   result_col75[30] <= result_col75[29];
   result_col75[31] <= result_col75[30];
   result_col75[32] <= result_col75[31];
   result_col75[33] <= result_col75[32];
   result_col75[34] <= result_col75[33];
   result_col75[35] <= result_col75[34];
   result_col75[36] <= result_col75[35];
   result_col75[37] <= result_col75[36];
   result_col75[38] <= result_col75[37];
   result_col75[39] <= result_col75[38];
   result_col75[40] <= result_col75[39];
   result_col75[41] <= result_col75[40];
   result_col75[42] <= result_col75[41];
   result_col75[43] <= result_col75[42];
   result_col75[44] <= result_col75[43];
   result_col75[45] <= result_col75[44];
   result_col75[46] <= result_col75[45];
   result_col75[47] <= result_col75[46];
   result_col75[48] <= result_col75[47];
   result_col75[49] <= result_col75[48];
   result_col75[50] <= result_col75[49];
   result_col75[51] <= result_col75[50];
   result_col75[52] <= result_col75[51];
   result_col75[53] <= result_col75[52];
   result_col75[54] <= result_col75[53];
   result_col75[55] <= result_col75[54];
   result_col75[56] <= result_col75[55];
   result_col75[57] <= result_col75[56];
   result_col75[58] <= result_col75[57];
   result_col75[59] <= result_col75[58];
   result_col75[60] <= result_col75[59];
   result_col75[61] <= result_col75[60];
   result_col75[62] <= result_col75[61];
   result_col75[63] <= result_col75[62];
   result_col75[64] <= result_col75[63];
   result_col75[65] <= result_col75[64];
   result_col75[66] <= result_col75[65];
   result_col75[67] <= result_col75[66];
   result_col75[68] <= result_col75[67];
   result_col75[69] <= result_col75[68];
   result_col75[70] <= result_col75[69];
   result_col75[71] <= result_col75[70];
   result_col75[72] <= result_col75[71];
   result_col75[73] <= result_col75[72];
   result_col75[74] <= result_col75[73];
   result_col75[75] <= result_col75[74];
   result_col75[76] <= result_col75[75];
   result_col75[77] <= result_col75[76];
   result_col75[78] <= result_col75[77];
   result_col75[79] <= result_col75[78];
   result_col75[80] <= result_col75[79];
   result_col75[81] <= result_col75[80];
   result_col75[82] <= result_col75[81];
   result_col75[83] <= result_col75[82];
   result_col75[84] <= result_col75[83];
   result_col75[85] <= result_col75[84];
   result_col75[86] <= result_col75[85];
   result_col75[87] <= result_col75[86];
   result_col75[88] <= result_col75[87];
   result_col75[89] <= result_col75[88];
   result_col75[90] <= result_col75[89];
   result_col75[91] <= result_col75[90];

   result_col76[1] <= data_out_4_76;
   result_col76[2] <= result_col76[1];
   result_col76[3] <= result_col76[2];
   result_col76[4] <= result_col76[3];
   result_col76[5] <= result_col76[4];
   result_col76[6] <= result_col76[5];
   result_col76[7] <= result_col76[6];
   result_col76[8] <= result_col76[7];
   result_col76[9] <= result_col76[8];
   result_col76[10] <= result_col76[9];
   result_col76[11] <= result_col76[10];
   result_col76[12] <= result_col76[11];
   result_col76[13] <= result_col76[12];
   result_col76[14] <= result_col76[13];
   result_col76[15] <= result_col76[14];
   result_col76[16] <= result_col76[15];
   result_col76[17] <= result_col76[16];
   result_col76[18] <= result_col76[17];
   result_col76[19] <= result_col76[18];
   result_col76[20] <= result_col76[19];
   result_col76[21] <= result_col76[20];
   result_col76[22] <= result_col76[21];
   result_col76[23] <= result_col76[22];
   result_col76[24] <= result_col76[23];
   result_col76[25] <= result_col76[24];
   result_col76[26] <= result_col76[25];
   result_col76[27] <= result_col76[26];
   result_col76[28] <= result_col76[27];
   result_col76[29] <= result_col76[28];
   result_col76[30] <= result_col76[29];
   result_col76[31] <= result_col76[30];
   result_col76[32] <= result_col76[31];
   result_col76[33] <= result_col76[32];
   result_col76[34] <= result_col76[33];
   result_col76[35] <= result_col76[34];
   result_col76[36] <= result_col76[35];
   result_col76[37] <= result_col76[36];
   result_col76[38] <= result_col76[37];
   result_col76[39] <= result_col76[38];
   result_col76[40] <= result_col76[39];
   result_col76[41] <= result_col76[40];
   result_col76[42] <= result_col76[41];
   result_col76[43] <= result_col76[42];
   result_col76[44] <= result_col76[43];
   result_col76[45] <= result_col76[44];
   result_col76[46] <= result_col76[45];
   result_col76[47] <= result_col76[46];
   result_col76[48] <= result_col76[47];
   result_col76[49] <= result_col76[48];
   result_col76[50] <= result_col76[49];
   result_col76[51] <= result_col76[50];
   result_col76[52] <= result_col76[51];
   result_col76[53] <= result_col76[52];
   result_col76[54] <= result_col76[53];
   result_col76[55] <= result_col76[54];
   result_col76[56] <= result_col76[55];
   result_col76[57] <= result_col76[56];
   result_col76[58] <= result_col76[57];
   result_col76[59] <= result_col76[58];
   result_col76[60] <= result_col76[59];
   result_col76[61] <= result_col76[60];
   result_col76[62] <= result_col76[61];
   result_col76[63] <= result_col76[62];
   result_col76[64] <= result_col76[63];
   result_col76[65] <= result_col76[64];
   result_col76[66] <= result_col76[65];
   result_col76[67] <= result_col76[66];
   result_col76[68] <= result_col76[67];
   result_col76[69] <= result_col76[68];
   result_col76[70] <= result_col76[69];
   result_col76[71] <= result_col76[70];
   result_col76[72] <= result_col76[71];
   result_col76[73] <= result_col76[72];
   result_col76[74] <= result_col76[73];
   result_col76[75] <= result_col76[74];
   result_col76[76] <= result_col76[75];
   result_col76[77] <= result_col76[76];
   result_col76[78] <= result_col76[77];
   result_col76[79] <= result_col76[78];
   result_col76[80] <= result_col76[79];
   result_col76[81] <= result_col76[80];
   result_col76[82] <= result_col76[81];
   result_col76[83] <= result_col76[82];
   result_col76[84] <= result_col76[83];
   result_col76[85] <= result_col76[84];
   result_col76[86] <= result_col76[85];
   result_col76[87] <= result_col76[86];
   result_col76[88] <= result_col76[87];
   result_col76[89] <= result_col76[88];
   result_col76[90] <= result_col76[89];

   result_col77[1] <= data_out_4_77;
   result_col77[2] <= result_col77[1];
   result_col77[3] <= result_col77[2];
   result_col77[4] <= result_col77[3];
   result_col77[5] <= result_col77[4];
   result_col77[6] <= result_col77[5];
   result_col77[7] <= result_col77[6];
   result_col77[8] <= result_col77[7];
   result_col77[9] <= result_col77[8];
   result_col77[10] <= result_col77[9];
   result_col77[11] <= result_col77[10];
   result_col77[12] <= result_col77[11];
   result_col77[13] <= result_col77[12];
   result_col77[14] <= result_col77[13];
   result_col77[15] <= result_col77[14];
   result_col77[16] <= result_col77[15];
   result_col77[17] <= result_col77[16];
   result_col77[18] <= result_col77[17];
   result_col77[19] <= result_col77[18];
   result_col77[20] <= result_col77[19];
   result_col77[21] <= result_col77[20];
   result_col77[22] <= result_col77[21];
   result_col77[23] <= result_col77[22];
   result_col77[24] <= result_col77[23];
   result_col77[25] <= result_col77[24];
   result_col77[26] <= result_col77[25];
   result_col77[27] <= result_col77[26];
   result_col77[28] <= result_col77[27];
   result_col77[29] <= result_col77[28];
   result_col77[30] <= result_col77[29];
   result_col77[31] <= result_col77[30];
   result_col77[32] <= result_col77[31];
   result_col77[33] <= result_col77[32];
   result_col77[34] <= result_col77[33];
   result_col77[35] <= result_col77[34];
   result_col77[36] <= result_col77[35];
   result_col77[37] <= result_col77[36];
   result_col77[38] <= result_col77[37];
   result_col77[39] <= result_col77[38];
   result_col77[40] <= result_col77[39];
   result_col77[41] <= result_col77[40];
   result_col77[42] <= result_col77[41];
   result_col77[43] <= result_col77[42];
   result_col77[44] <= result_col77[43];
   result_col77[45] <= result_col77[44];
   result_col77[46] <= result_col77[45];
   result_col77[47] <= result_col77[46];
   result_col77[48] <= result_col77[47];
   result_col77[49] <= result_col77[48];
   result_col77[50] <= result_col77[49];
   result_col77[51] <= result_col77[50];
   result_col77[52] <= result_col77[51];
   result_col77[53] <= result_col77[52];
   result_col77[54] <= result_col77[53];
   result_col77[55] <= result_col77[54];
   result_col77[56] <= result_col77[55];
   result_col77[57] <= result_col77[56];
   result_col77[58] <= result_col77[57];
   result_col77[59] <= result_col77[58];
   result_col77[60] <= result_col77[59];
   result_col77[61] <= result_col77[60];
   result_col77[62] <= result_col77[61];
   result_col77[63] <= result_col77[62];
   result_col77[64] <= result_col77[63];
   result_col77[65] <= result_col77[64];
   result_col77[66] <= result_col77[65];
   result_col77[67] <= result_col77[66];
   result_col77[68] <= result_col77[67];
   result_col77[69] <= result_col77[68];
   result_col77[70] <= result_col77[69];
   result_col77[71] <= result_col77[70];
   result_col77[72] <= result_col77[71];
   result_col77[73] <= result_col77[72];
   result_col77[74] <= result_col77[73];
   result_col77[75] <= result_col77[74];
   result_col77[76] <= result_col77[75];
   result_col77[77] <= result_col77[76];
   result_col77[78] <= result_col77[77];
   result_col77[79] <= result_col77[78];
   result_col77[80] <= result_col77[79];
   result_col77[81] <= result_col77[80];
   result_col77[82] <= result_col77[81];
   result_col77[83] <= result_col77[82];
   result_col77[84] <= result_col77[83];
   result_col77[85] <= result_col77[84];
   result_col77[86] <= result_col77[85];
   result_col77[87] <= result_col77[86];
   result_col77[88] <= result_col77[87];
   result_col77[89] <= result_col77[88];

   result_col78[1] <= data_out_4_78;
   result_col78[2] <= result_col78[1];
   result_col78[3] <= result_col78[2];
   result_col78[4] <= result_col78[3];
   result_col78[5] <= result_col78[4];
   result_col78[6] <= result_col78[5];
   result_col78[7] <= result_col78[6];
   result_col78[8] <= result_col78[7];
   result_col78[9] <= result_col78[8];
   result_col78[10] <= result_col78[9];
   result_col78[11] <= result_col78[10];
   result_col78[12] <= result_col78[11];
   result_col78[13] <= result_col78[12];
   result_col78[14] <= result_col78[13];
   result_col78[15] <= result_col78[14];
   result_col78[16] <= result_col78[15];
   result_col78[17] <= result_col78[16];
   result_col78[18] <= result_col78[17];
   result_col78[19] <= result_col78[18];
   result_col78[20] <= result_col78[19];
   result_col78[21] <= result_col78[20];
   result_col78[22] <= result_col78[21];
   result_col78[23] <= result_col78[22];
   result_col78[24] <= result_col78[23];
   result_col78[25] <= result_col78[24];
   result_col78[26] <= result_col78[25];
   result_col78[27] <= result_col78[26];
   result_col78[28] <= result_col78[27];
   result_col78[29] <= result_col78[28];
   result_col78[30] <= result_col78[29];
   result_col78[31] <= result_col78[30];
   result_col78[32] <= result_col78[31];
   result_col78[33] <= result_col78[32];
   result_col78[34] <= result_col78[33];
   result_col78[35] <= result_col78[34];
   result_col78[36] <= result_col78[35];
   result_col78[37] <= result_col78[36];
   result_col78[38] <= result_col78[37];
   result_col78[39] <= result_col78[38];
   result_col78[40] <= result_col78[39];
   result_col78[41] <= result_col78[40];
   result_col78[42] <= result_col78[41];
   result_col78[43] <= result_col78[42];
   result_col78[44] <= result_col78[43];
   result_col78[45] <= result_col78[44];
   result_col78[46] <= result_col78[45];
   result_col78[47] <= result_col78[46];
   result_col78[48] <= result_col78[47];
   result_col78[49] <= result_col78[48];
   result_col78[50] <= result_col78[49];
   result_col78[51] <= result_col78[50];
   result_col78[52] <= result_col78[51];
   result_col78[53] <= result_col78[52];
   result_col78[54] <= result_col78[53];
   result_col78[55] <= result_col78[54];
   result_col78[56] <= result_col78[55];
   result_col78[57] <= result_col78[56];
   result_col78[58] <= result_col78[57];
   result_col78[59] <= result_col78[58];
   result_col78[60] <= result_col78[59];
   result_col78[61] <= result_col78[60];
   result_col78[62] <= result_col78[61];
   result_col78[63] <= result_col78[62];
   result_col78[64] <= result_col78[63];
   result_col78[65] <= result_col78[64];
   result_col78[66] <= result_col78[65];
   result_col78[67] <= result_col78[66];
   result_col78[68] <= result_col78[67];
   result_col78[69] <= result_col78[68];
   result_col78[70] <= result_col78[69];
   result_col78[71] <= result_col78[70];
   result_col78[72] <= result_col78[71];
   result_col78[73] <= result_col78[72];
   result_col78[74] <= result_col78[73];
   result_col78[75] <= result_col78[74];
   result_col78[76] <= result_col78[75];
   result_col78[77] <= result_col78[76];
   result_col78[78] <= result_col78[77];
   result_col78[79] <= result_col78[78];
   result_col78[80] <= result_col78[79];
   result_col78[81] <= result_col78[80];
   result_col78[82] <= result_col78[81];
   result_col78[83] <= result_col78[82];
   result_col78[84] <= result_col78[83];
   result_col78[85] <= result_col78[84];
   result_col78[86] <= result_col78[85];
   result_col78[87] <= result_col78[86];
   result_col78[88] <= result_col78[87];

   result_col79[1] <= data_out_4_79;
   result_col79[2] <= result_col79[1];
   result_col79[3] <= result_col79[2];
   result_col79[4] <= result_col79[3];
   result_col79[5] <= result_col79[4];
   result_col79[6] <= result_col79[5];
   result_col79[7] <= result_col79[6];
   result_col79[8] <= result_col79[7];
   result_col79[9] <= result_col79[8];
   result_col79[10] <= result_col79[9];
   result_col79[11] <= result_col79[10];
   result_col79[12] <= result_col79[11];
   result_col79[13] <= result_col79[12];
   result_col79[14] <= result_col79[13];
   result_col79[15] <= result_col79[14];
   result_col79[16] <= result_col79[15];
   result_col79[17] <= result_col79[16];
   result_col79[18] <= result_col79[17];
   result_col79[19] <= result_col79[18];
   result_col79[20] <= result_col79[19];
   result_col79[21] <= result_col79[20];
   result_col79[22] <= result_col79[21];
   result_col79[23] <= result_col79[22];
   result_col79[24] <= result_col79[23];
   result_col79[25] <= result_col79[24];
   result_col79[26] <= result_col79[25];
   result_col79[27] <= result_col79[26];
   result_col79[28] <= result_col79[27];
   result_col79[29] <= result_col79[28];
   result_col79[30] <= result_col79[29];
   result_col79[31] <= result_col79[30];
   result_col79[32] <= result_col79[31];
   result_col79[33] <= result_col79[32];
   result_col79[34] <= result_col79[33];
   result_col79[35] <= result_col79[34];
   result_col79[36] <= result_col79[35];
   result_col79[37] <= result_col79[36];
   result_col79[38] <= result_col79[37];
   result_col79[39] <= result_col79[38];
   result_col79[40] <= result_col79[39];
   result_col79[41] <= result_col79[40];
   result_col79[42] <= result_col79[41];
   result_col79[43] <= result_col79[42];
   result_col79[44] <= result_col79[43];
   result_col79[45] <= result_col79[44];
   result_col79[46] <= result_col79[45];
   result_col79[47] <= result_col79[46];
   result_col79[48] <= result_col79[47];
   result_col79[49] <= result_col79[48];
   result_col79[50] <= result_col79[49];
   result_col79[51] <= result_col79[50];
   result_col79[52] <= result_col79[51];
   result_col79[53] <= result_col79[52];
   result_col79[54] <= result_col79[53];
   result_col79[55] <= result_col79[54];
   result_col79[56] <= result_col79[55];
   result_col79[57] <= result_col79[56];
   result_col79[58] <= result_col79[57];
   result_col79[59] <= result_col79[58];
   result_col79[60] <= result_col79[59];
   result_col79[61] <= result_col79[60];
   result_col79[62] <= result_col79[61];
   result_col79[63] <= result_col79[62];
   result_col79[64] <= result_col79[63];
   result_col79[65] <= result_col79[64];
   result_col79[66] <= result_col79[65];
   result_col79[67] <= result_col79[66];
   result_col79[68] <= result_col79[67];
   result_col79[69] <= result_col79[68];
   result_col79[70] <= result_col79[69];
   result_col79[71] <= result_col79[70];
   result_col79[72] <= result_col79[71];
   result_col79[73] <= result_col79[72];
   result_col79[74] <= result_col79[73];
   result_col79[75] <= result_col79[74];
   result_col79[76] <= result_col79[75];
   result_col79[77] <= result_col79[76];
   result_col79[78] <= result_col79[77];
   result_col79[79] <= result_col79[78];
   result_col79[80] <= result_col79[79];
   result_col79[81] <= result_col79[80];
   result_col79[82] <= result_col79[81];
   result_col79[83] <= result_col79[82];
   result_col79[84] <= result_col79[83];
   result_col79[85] <= result_col79[84];
   result_col79[86] <= result_col79[85];
   result_col79[87] <= result_col79[86];

   result_col80[1] <= data_out_4_80;
   result_col80[2] <= result_col80[1];
   result_col80[3] <= result_col80[2];
   result_col80[4] <= result_col80[3];
   result_col80[5] <= result_col80[4];
   result_col80[6] <= result_col80[5];
   result_col80[7] <= result_col80[6];
   result_col80[8] <= result_col80[7];
   result_col80[9] <= result_col80[8];
   result_col80[10] <= result_col80[9];
   result_col80[11] <= result_col80[10];
   result_col80[12] <= result_col80[11];
   result_col80[13] <= result_col80[12];
   result_col80[14] <= result_col80[13];
   result_col80[15] <= result_col80[14];
   result_col80[16] <= result_col80[15];
   result_col80[17] <= result_col80[16];
   result_col80[18] <= result_col80[17];
   result_col80[19] <= result_col80[18];
   result_col80[20] <= result_col80[19];
   result_col80[21] <= result_col80[20];
   result_col80[22] <= result_col80[21];
   result_col80[23] <= result_col80[22];
   result_col80[24] <= result_col80[23];
   result_col80[25] <= result_col80[24];
   result_col80[26] <= result_col80[25];
   result_col80[27] <= result_col80[26];
   result_col80[28] <= result_col80[27];
   result_col80[29] <= result_col80[28];
   result_col80[30] <= result_col80[29];
   result_col80[31] <= result_col80[30];
   result_col80[32] <= result_col80[31];
   result_col80[33] <= result_col80[32];
   result_col80[34] <= result_col80[33];
   result_col80[35] <= result_col80[34];
   result_col80[36] <= result_col80[35];
   result_col80[37] <= result_col80[36];
   result_col80[38] <= result_col80[37];
   result_col80[39] <= result_col80[38];
   result_col80[40] <= result_col80[39];
   result_col80[41] <= result_col80[40];
   result_col80[42] <= result_col80[41];
   result_col80[43] <= result_col80[42];
   result_col80[44] <= result_col80[43];
   result_col80[45] <= result_col80[44];
   result_col80[46] <= result_col80[45];
   result_col80[47] <= result_col80[46];
   result_col80[48] <= result_col80[47];
   result_col80[49] <= result_col80[48];
   result_col80[50] <= result_col80[49];
   result_col80[51] <= result_col80[50];
   result_col80[52] <= result_col80[51];
   result_col80[53] <= result_col80[52];
   result_col80[54] <= result_col80[53];
   result_col80[55] <= result_col80[54];
   result_col80[56] <= result_col80[55];
   result_col80[57] <= result_col80[56];
   result_col80[58] <= result_col80[57];
   result_col80[59] <= result_col80[58];
   result_col80[60] <= result_col80[59];
   result_col80[61] <= result_col80[60];
   result_col80[62] <= result_col80[61];
   result_col80[63] <= result_col80[62];
   result_col80[64] <= result_col80[63];
   result_col80[65] <= result_col80[64];
   result_col80[66] <= result_col80[65];
   result_col80[67] <= result_col80[66];
   result_col80[68] <= result_col80[67];
   result_col80[69] <= result_col80[68];
   result_col80[70] <= result_col80[69];
   result_col80[71] <= result_col80[70];
   result_col80[72] <= result_col80[71];
   result_col80[73] <= result_col80[72];
   result_col80[74] <= result_col80[73];
   result_col80[75] <= result_col80[74];
   result_col80[76] <= result_col80[75];
   result_col80[77] <= result_col80[76];
   result_col80[78] <= result_col80[77];
   result_col80[79] <= result_col80[78];
   result_col80[80] <= result_col80[79];
   result_col80[81] <= result_col80[80];
   result_col80[82] <= result_col80[81];
   result_col80[83] <= result_col80[82];
   result_col80[84] <= result_col80[83];
   result_col80[85] <= result_col80[84];
   result_col80[86] <= result_col80[85];

   result_col81[1] <= data_out_4_81;
   result_col81[2] <= result_col81[1];
   result_col81[3] <= result_col81[2];
   result_col81[4] <= result_col81[3];
   result_col81[5] <= result_col81[4];
   result_col81[6] <= result_col81[5];
   result_col81[7] <= result_col81[6];
   result_col81[8] <= result_col81[7];
   result_col81[9] <= result_col81[8];
   result_col81[10] <= result_col81[9];
   result_col81[11] <= result_col81[10];
   result_col81[12] <= result_col81[11];
   result_col81[13] <= result_col81[12];
   result_col81[14] <= result_col81[13];
   result_col81[15] <= result_col81[14];
   result_col81[16] <= result_col81[15];
   result_col81[17] <= result_col81[16];
   result_col81[18] <= result_col81[17];
   result_col81[19] <= result_col81[18];
   result_col81[20] <= result_col81[19];
   result_col81[21] <= result_col81[20];
   result_col81[22] <= result_col81[21];
   result_col81[23] <= result_col81[22];
   result_col81[24] <= result_col81[23];
   result_col81[25] <= result_col81[24];
   result_col81[26] <= result_col81[25];
   result_col81[27] <= result_col81[26];
   result_col81[28] <= result_col81[27];
   result_col81[29] <= result_col81[28];
   result_col81[30] <= result_col81[29];
   result_col81[31] <= result_col81[30];
   result_col81[32] <= result_col81[31];
   result_col81[33] <= result_col81[32];
   result_col81[34] <= result_col81[33];
   result_col81[35] <= result_col81[34];
   result_col81[36] <= result_col81[35];
   result_col81[37] <= result_col81[36];
   result_col81[38] <= result_col81[37];
   result_col81[39] <= result_col81[38];
   result_col81[40] <= result_col81[39];
   result_col81[41] <= result_col81[40];
   result_col81[42] <= result_col81[41];
   result_col81[43] <= result_col81[42];
   result_col81[44] <= result_col81[43];
   result_col81[45] <= result_col81[44];
   result_col81[46] <= result_col81[45];
   result_col81[47] <= result_col81[46];
   result_col81[48] <= result_col81[47];
   result_col81[49] <= result_col81[48];
   result_col81[50] <= result_col81[49];
   result_col81[51] <= result_col81[50];
   result_col81[52] <= result_col81[51];
   result_col81[53] <= result_col81[52];
   result_col81[54] <= result_col81[53];
   result_col81[55] <= result_col81[54];
   result_col81[56] <= result_col81[55];
   result_col81[57] <= result_col81[56];
   result_col81[58] <= result_col81[57];
   result_col81[59] <= result_col81[58];
   result_col81[60] <= result_col81[59];
   result_col81[61] <= result_col81[60];
   result_col81[62] <= result_col81[61];
   result_col81[63] <= result_col81[62];
   result_col81[64] <= result_col81[63];
   result_col81[65] <= result_col81[64];
   result_col81[66] <= result_col81[65];
   result_col81[67] <= result_col81[66];
   result_col81[68] <= result_col81[67];
   result_col81[69] <= result_col81[68];
   result_col81[70] <= result_col81[69];
   result_col81[71] <= result_col81[70];
   result_col81[72] <= result_col81[71];
   result_col81[73] <= result_col81[72];
   result_col81[74] <= result_col81[73];
   result_col81[75] <= result_col81[74];
   result_col81[76] <= result_col81[75];
   result_col81[77] <= result_col81[76];
   result_col81[78] <= result_col81[77];
   result_col81[79] <= result_col81[78];
   result_col81[80] <= result_col81[79];
   result_col81[81] <= result_col81[80];
   result_col81[82] <= result_col81[81];
   result_col81[83] <= result_col81[82];
   result_col81[84] <= result_col81[83];
   result_col81[85] <= result_col81[84];

   result_col82[1] <= data_out_4_82;
   result_col82[2] <= result_col82[1];
   result_col82[3] <= result_col82[2];
   result_col82[4] <= result_col82[3];
   result_col82[5] <= result_col82[4];
   result_col82[6] <= result_col82[5];
   result_col82[7] <= result_col82[6];
   result_col82[8] <= result_col82[7];
   result_col82[9] <= result_col82[8];
   result_col82[10] <= result_col82[9];
   result_col82[11] <= result_col82[10];
   result_col82[12] <= result_col82[11];
   result_col82[13] <= result_col82[12];
   result_col82[14] <= result_col82[13];
   result_col82[15] <= result_col82[14];
   result_col82[16] <= result_col82[15];
   result_col82[17] <= result_col82[16];
   result_col82[18] <= result_col82[17];
   result_col82[19] <= result_col82[18];
   result_col82[20] <= result_col82[19];
   result_col82[21] <= result_col82[20];
   result_col82[22] <= result_col82[21];
   result_col82[23] <= result_col82[22];
   result_col82[24] <= result_col82[23];
   result_col82[25] <= result_col82[24];
   result_col82[26] <= result_col82[25];
   result_col82[27] <= result_col82[26];
   result_col82[28] <= result_col82[27];
   result_col82[29] <= result_col82[28];
   result_col82[30] <= result_col82[29];
   result_col82[31] <= result_col82[30];
   result_col82[32] <= result_col82[31];
   result_col82[33] <= result_col82[32];
   result_col82[34] <= result_col82[33];
   result_col82[35] <= result_col82[34];
   result_col82[36] <= result_col82[35];
   result_col82[37] <= result_col82[36];
   result_col82[38] <= result_col82[37];
   result_col82[39] <= result_col82[38];
   result_col82[40] <= result_col82[39];
   result_col82[41] <= result_col82[40];
   result_col82[42] <= result_col82[41];
   result_col82[43] <= result_col82[42];
   result_col82[44] <= result_col82[43];
   result_col82[45] <= result_col82[44];
   result_col82[46] <= result_col82[45];
   result_col82[47] <= result_col82[46];
   result_col82[48] <= result_col82[47];
   result_col82[49] <= result_col82[48];
   result_col82[50] <= result_col82[49];
   result_col82[51] <= result_col82[50];
   result_col82[52] <= result_col82[51];
   result_col82[53] <= result_col82[52];
   result_col82[54] <= result_col82[53];
   result_col82[55] <= result_col82[54];
   result_col82[56] <= result_col82[55];
   result_col82[57] <= result_col82[56];
   result_col82[58] <= result_col82[57];
   result_col82[59] <= result_col82[58];
   result_col82[60] <= result_col82[59];
   result_col82[61] <= result_col82[60];
   result_col82[62] <= result_col82[61];
   result_col82[63] <= result_col82[62];
   result_col82[64] <= result_col82[63];
   result_col82[65] <= result_col82[64];
   result_col82[66] <= result_col82[65];
   result_col82[67] <= result_col82[66];
   result_col82[68] <= result_col82[67];
   result_col82[69] <= result_col82[68];
   result_col82[70] <= result_col82[69];
   result_col82[71] <= result_col82[70];
   result_col82[72] <= result_col82[71];
   result_col82[73] <= result_col82[72];
   result_col82[74] <= result_col82[73];
   result_col82[75] <= result_col82[74];
   result_col82[76] <= result_col82[75];
   result_col82[77] <= result_col82[76];
   result_col82[78] <= result_col82[77];
   result_col82[79] <= result_col82[78];
   result_col82[80] <= result_col82[79];
   result_col82[81] <= result_col82[80];
   result_col82[82] <= result_col82[81];
   result_col82[83] <= result_col82[82];
   result_col82[84] <= result_col82[83];

   result_col83[1] <= data_out_4_83;
   result_col83[2] <= result_col83[1];
   result_col83[3] <= result_col83[2];
   result_col83[4] <= result_col83[3];
   result_col83[5] <= result_col83[4];
   result_col83[6] <= result_col83[5];
   result_col83[7] <= result_col83[6];
   result_col83[8] <= result_col83[7];
   result_col83[9] <= result_col83[8];
   result_col83[10] <= result_col83[9];
   result_col83[11] <= result_col83[10];
   result_col83[12] <= result_col83[11];
   result_col83[13] <= result_col83[12];
   result_col83[14] <= result_col83[13];
   result_col83[15] <= result_col83[14];
   result_col83[16] <= result_col83[15];
   result_col83[17] <= result_col83[16];
   result_col83[18] <= result_col83[17];
   result_col83[19] <= result_col83[18];
   result_col83[20] <= result_col83[19];
   result_col83[21] <= result_col83[20];
   result_col83[22] <= result_col83[21];
   result_col83[23] <= result_col83[22];
   result_col83[24] <= result_col83[23];
   result_col83[25] <= result_col83[24];
   result_col83[26] <= result_col83[25];
   result_col83[27] <= result_col83[26];
   result_col83[28] <= result_col83[27];
   result_col83[29] <= result_col83[28];
   result_col83[30] <= result_col83[29];
   result_col83[31] <= result_col83[30];
   result_col83[32] <= result_col83[31];
   result_col83[33] <= result_col83[32];
   result_col83[34] <= result_col83[33];
   result_col83[35] <= result_col83[34];
   result_col83[36] <= result_col83[35];
   result_col83[37] <= result_col83[36];
   result_col83[38] <= result_col83[37];
   result_col83[39] <= result_col83[38];
   result_col83[40] <= result_col83[39];
   result_col83[41] <= result_col83[40];
   result_col83[42] <= result_col83[41];
   result_col83[43] <= result_col83[42];
   result_col83[44] <= result_col83[43];
   result_col83[45] <= result_col83[44];
   result_col83[46] <= result_col83[45];
   result_col83[47] <= result_col83[46];
   result_col83[48] <= result_col83[47];
   result_col83[49] <= result_col83[48];
   result_col83[50] <= result_col83[49];
   result_col83[51] <= result_col83[50];
   result_col83[52] <= result_col83[51];
   result_col83[53] <= result_col83[52];
   result_col83[54] <= result_col83[53];
   result_col83[55] <= result_col83[54];
   result_col83[56] <= result_col83[55];
   result_col83[57] <= result_col83[56];
   result_col83[58] <= result_col83[57];
   result_col83[59] <= result_col83[58];
   result_col83[60] <= result_col83[59];
   result_col83[61] <= result_col83[60];
   result_col83[62] <= result_col83[61];
   result_col83[63] <= result_col83[62];
   result_col83[64] <= result_col83[63];
   result_col83[65] <= result_col83[64];
   result_col83[66] <= result_col83[65];
   result_col83[67] <= result_col83[66];
   result_col83[68] <= result_col83[67];
   result_col83[69] <= result_col83[68];
   result_col83[70] <= result_col83[69];
   result_col83[71] <= result_col83[70];
   result_col83[72] <= result_col83[71];
   result_col83[73] <= result_col83[72];
   result_col83[74] <= result_col83[73];
   result_col83[75] <= result_col83[74];
   result_col83[76] <= result_col83[75];
   result_col83[77] <= result_col83[76];
   result_col83[78] <= result_col83[77];
   result_col83[79] <= result_col83[78];
   result_col83[80] <= result_col83[79];
   result_col83[81] <= result_col83[80];
   result_col83[82] <= result_col83[81];
   result_col83[83] <= result_col83[82];

   result_col84[1] <= data_out_4_84;
   result_col84[2] <= result_col84[1];
   result_col84[3] <= result_col84[2];
   result_col84[4] <= result_col84[3];
   result_col84[5] <= result_col84[4];
   result_col84[6] <= result_col84[5];
   result_col84[7] <= result_col84[6];
   result_col84[8] <= result_col84[7];
   result_col84[9] <= result_col84[8];
   result_col84[10] <= result_col84[9];
   result_col84[11] <= result_col84[10];
   result_col84[12] <= result_col84[11];
   result_col84[13] <= result_col84[12];
   result_col84[14] <= result_col84[13];
   result_col84[15] <= result_col84[14];
   result_col84[16] <= result_col84[15];
   result_col84[17] <= result_col84[16];
   result_col84[18] <= result_col84[17];
   result_col84[19] <= result_col84[18];
   result_col84[20] <= result_col84[19];
   result_col84[21] <= result_col84[20];
   result_col84[22] <= result_col84[21];
   result_col84[23] <= result_col84[22];
   result_col84[24] <= result_col84[23];
   result_col84[25] <= result_col84[24];
   result_col84[26] <= result_col84[25];
   result_col84[27] <= result_col84[26];
   result_col84[28] <= result_col84[27];
   result_col84[29] <= result_col84[28];
   result_col84[30] <= result_col84[29];
   result_col84[31] <= result_col84[30];
   result_col84[32] <= result_col84[31];
   result_col84[33] <= result_col84[32];
   result_col84[34] <= result_col84[33];
   result_col84[35] <= result_col84[34];
   result_col84[36] <= result_col84[35];
   result_col84[37] <= result_col84[36];
   result_col84[38] <= result_col84[37];
   result_col84[39] <= result_col84[38];
   result_col84[40] <= result_col84[39];
   result_col84[41] <= result_col84[40];
   result_col84[42] <= result_col84[41];
   result_col84[43] <= result_col84[42];
   result_col84[44] <= result_col84[43];
   result_col84[45] <= result_col84[44];
   result_col84[46] <= result_col84[45];
   result_col84[47] <= result_col84[46];
   result_col84[48] <= result_col84[47];
   result_col84[49] <= result_col84[48];
   result_col84[50] <= result_col84[49];
   result_col84[51] <= result_col84[50];
   result_col84[52] <= result_col84[51];
   result_col84[53] <= result_col84[52];
   result_col84[54] <= result_col84[53];
   result_col84[55] <= result_col84[54];
   result_col84[56] <= result_col84[55];
   result_col84[57] <= result_col84[56];
   result_col84[58] <= result_col84[57];
   result_col84[59] <= result_col84[58];
   result_col84[60] <= result_col84[59];
   result_col84[61] <= result_col84[60];
   result_col84[62] <= result_col84[61];
   result_col84[63] <= result_col84[62];
   result_col84[64] <= result_col84[63];
   result_col84[65] <= result_col84[64];
   result_col84[66] <= result_col84[65];
   result_col84[67] <= result_col84[66];
   result_col84[68] <= result_col84[67];
   result_col84[69] <= result_col84[68];
   result_col84[70] <= result_col84[69];
   result_col84[71] <= result_col84[70];
   result_col84[72] <= result_col84[71];
   result_col84[73] <= result_col84[72];
   result_col84[74] <= result_col84[73];
   result_col84[75] <= result_col84[74];
   result_col84[76] <= result_col84[75];
   result_col84[77] <= result_col84[76];
   result_col84[78] <= result_col84[77];
   result_col84[79] <= result_col84[78];
   result_col84[80] <= result_col84[79];
   result_col84[81] <= result_col84[80];
   result_col84[82] <= result_col84[81];

   result_col85[1] <= data_out_4_85;
   result_col85[2] <= result_col85[1];
   result_col85[3] <= result_col85[2];
   result_col85[4] <= result_col85[3];
   result_col85[5] <= result_col85[4];
   result_col85[6] <= result_col85[5];
   result_col85[7] <= result_col85[6];
   result_col85[8] <= result_col85[7];
   result_col85[9] <= result_col85[8];
   result_col85[10] <= result_col85[9];
   result_col85[11] <= result_col85[10];
   result_col85[12] <= result_col85[11];
   result_col85[13] <= result_col85[12];
   result_col85[14] <= result_col85[13];
   result_col85[15] <= result_col85[14];
   result_col85[16] <= result_col85[15];
   result_col85[17] <= result_col85[16];
   result_col85[18] <= result_col85[17];
   result_col85[19] <= result_col85[18];
   result_col85[20] <= result_col85[19];
   result_col85[21] <= result_col85[20];
   result_col85[22] <= result_col85[21];
   result_col85[23] <= result_col85[22];
   result_col85[24] <= result_col85[23];
   result_col85[25] <= result_col85[24];
   result_col85[26] <= result_col85[25];
   result_col85[27] <= result_col85[26];
   result_col85[28] <= result_col85[27];
   result_col85[29] <= result_col85[28];
   result_col85[30] <= result_col85[29];
   result_col85[31] <= result_col85[30];
   result_col85[32] <= result_col85[31];
   result_col85[33] <= result_col85[32];
   result_col85[34] <= result_col85[33];
   result_col85[35] <= result_col85[34];
   result_col85[36] <= result_col85[35];
   result_col85[37] <= result_col85[36];
   result_col85[38] <= result_col85[37];
   result_col85[39] <= result_col85[38];
   result_col85[40] <= result_col85[39];
   result_col85[41] <= result_col85[40];
   result_col85[42] <= result_col85[41];
   result_col85[43] <= result_col85[42];
   result_col85[44] <= result_col85[43];
   result_col85[45] <= result_col85[44];
   result_col85[46] <= result_col85[45];
   result_col85[47] <= result_col85[46];
   result_col85[48] <= result_col85[47];
   result_col85[49] <= result_col85[48];
   result_col85[50] <= result_col85[49];
   result_col85[51] <= result_col85[50];
   result_col85[52] <= result_col85[51];
   result_col85[53] <= result_col85[52];
   result_col85[54] <= result_col85[53];
   result_col85[55] <= result_col85[54];
   result_col85[56] <= result_col85[55];
   result_col85[57] <= result_col85[56];
   result_col85[58] <= result_col85[57];
   result_col85[59] <= result_col85[58];
   result_col85[60] <= result_col85[59];
   result_col85[61] <= result_col85[60];
   result_col85[62] <= result_col85[61];
   result_col85[63] <= result_col85[62];
   result_col85[64] <= result_col85[63];
   result_col85[65] <= result_col85[64];
   result_col85[66] <= result_col85[65];
   result_col85[67] <= result_col85[66];
   result_col85[68] <= result_col85[67];
   result_col85[69] <= result_col85[68];
   result_col85[70] <= result_col85[69];
   result_col85[71] <= result_col85[70];
   result_col85[72] <= result_col85[71];
   result_col85[73] <= result_col85[72];
   result_col85[74] <= result_col85[73];
   result_col85[75] <= result_col85[74];
   result_col85[76] <= result_col85[75];
   result_col85[77] <= result_col85[76];
   result_col85[78] <= result_col85[77];
   result_col85[79] <= result_col85[78];
   result_col85[80] <= result_col85[79];
   result_col85[81] <= result_col85[80];

   result_col86[1] <= data_out_4_86;
   result_col86[2] <= result_col86[1];
   result_col86[3] <= result_col86[2];
   result_col86[4] <= result_col86[3];
   result_col86[5] <= result_col86[4];
   result_col86[6] <= result_col86[5];
   result_col86[7] <= result_col86[6];
   result_col86[8] <= result_col86[7];
   result_col86[9] <= result_col86[8];
   result_col86[10] <= result_col86[9];
   result_col86[11] <= result_col86[10];
   result_col86[12] <= result_col86[11];
   result_col86[13] <= result_col86[12];
   result_col86[14] <= result_col86[13];
   result_col86[15] <= result_col86[14];
   result_col86[16] <= result_col86[15];
   result_col86[17] <= result_col86[16];
   result_col86[18] <= result_col86[17];
   result_col86[19] <= result_col86[18];
   result_col86[20] <= result_col86[19];
   result_col86[21] <= result_col86[20];
   result_col86[22] <= result_col86[21];
   result_col86[23] <= result_col86[22];
   result_col86[24] <= result_col86[23];
   result_col86[25] <= result_col86[24];
   result_col86[26] <= result_col86[25];
   result_col86[27] <= result_col86[26];
   result_col86[28] <= result_col86[27];
   result_col86[29] <= result_col86[28];
   result_col86[30] <= result_col86[29];
   result_col86[31] <= result_col86[30];
   result_col86[32] <= result_col86[31];
   result_col86[33] <= result_col86[32];
   result_col86[34] <= result_col86[33];
   result_col86[35] <= result_col86[34];
   result_col86[36] <= result_col86[35];
   result_col86[37] <= result_col86[36];
   result_col86[38] <= result_col86[37];
   result_col86[39] <= result_col86[38];
   result_col86[40] <= result_col86[39];
   result_col86[41] <= result_col86[40];
   result_col86[42] <= result_col86[41];
   result_col86[43] <= result_col86[42];
   result_col86[44] <= result_col86[43];
   result_col86[45] <= result_col86[44];
   result_col86[46] <= result_col86[45];
   result_col86[47] <= result_col86[46];
   result_col86[48] <= result_col86[47];
   result_col86[49] <= result_col86[48];
   result_col86[50] <= result_col86[49];
   result_col86[51] <= result_col86[50];
   result_col86[52] <= result_col86[51];
   result_col86[53] <= result_col86[52];
   result_col86[54] <= result_col86[53];
   result_col86[55] <= result_col86[54];
   result_col86[56] <= result_col86[55];
   result_col86[57] <= result_col86[56];
   result_col86[58] <= result_col86[57];
   result_col86[59] <= result_col86[58];
   result_col86[60] <= result_col86[59];
   result_col86[61] <= result_col86[60];
   result_col86[62] <= result_col86[61];
   result_col86[63] <= result_col86[62];
   result_col86[64] <= result_col86[63];
   result_col86[65] <= result_col86[64];
   result_col86[66] <= result_col86[65];
   result_col86[67] <= result_col86[66];
   result_col86[68] <= result_col86[67];
   result_col86[69] <= result_col86[68];
   result_col86[70] <= result_col86[69];
   result_col86[71] <= result_col86[70];
   result_col86[72] <= result_col86[71];
   result_col86[73] <= result_col86[72];
   result_col86[74] <= result_col86[73];
   result_col86[75] <= result_col86[74];
   result_col86[76] <= result_col86[75];
   result_col86[77] <= result_col86[76];
   result_col86[78] <= result_col86[77];
   result_col86[79] <= result_col86[78];
   result_col86[80] <= result_col86[79];

   result_col87[1] <= data_out_4_87;
   result_col87[2] <= result_col87[1];
   result_col87[3] <= result_col87[2];
   result_col87[4] <= result_col87[3];
   result_col87[5] <= result_col87[4];
   result_col87[6] <= result_col87[5];
   result_col87[7] <= result_col87[6];
   result_col87[8] <= result_col87[7];
   result_col87[9] <= result_col87[8];
   result_col87[10] <= result_col87[9];
   result_col87[11] <= result_col87[10];
   result_col87[12] <= result_col87[11];
   result_col87[13] <= result_col87[12];
   result_col87[14] <= result_col87[13];
   result_col87[15] <= result_col87[14];
   result_col87[16] <= result_col87[15];
   result_col87[17] <= result_col87[16];
   result_col87[18] <= result_col87[17];
   result_col87[19] <= result_col87[18];
   result_col87[20] <= result_col87[19];
   result_col87[21] <= result_col87[20];
   result_col87[22] <= result_col87[21];
   result_col87[23] <= result_col87[22];
   result_col87[24] <= result_col87[23];
   result_col87[25] <= result_col87[24];
   result_col87[26] <= result_col87[25];
   result_col87[27] <= result_col87[26];
   result_col87[28] <= result_col87[27];
   result_col87[29] <= result_col87[28];
   result_col87[30] <= result_col87[29];
   result_col87[31] <= result_col87[30];
   result_col87[32] <= result_col87[31];
   result_col87[33] <= result_col87[32];
   result_col87[34] <= result_col87[33];
   result_col87[35] <= result_col87[34];
   result_col87[36] <= result_col87[35];
   result_col87[37] <= result_col87[36];
   result_col87[38] <= result_col87[37];
   result_col87[39] <= result_col87[38];
   result_col87[40] <= result_col87[39];
   result_col87[41] <= result_col87[40];
   result_col87[42] <= result_col87[41];
   result_col87[43] <= result_col87[42];
   result_col87[44] <= result_col87[43];
   result_col87[45] <= result_col87[44];
   result_col87[46] <= result_col87[45];
   result_col87[47] <= result_col87[46];
   result_col87[48] <= result_col87[47];
   result_col87[49] <= result_col87[48];
   result_col87[50] <= result_col87[49];
   result_col87[51] <= result_col87[50];
   result_col87[52] <= result_col87[51];
   result_col87[53] <= result_col87[52];
   result_col87[54] <= result_col87[53];
   result_col87[55] <= result_col87[54];
   result_col87[56] <= result_col87[55];
   result_col87[57] <= result_col87[56];
   result_col87[58] <= result_col87[57];
   result_col87[59] <= result_col87[58];
   result_col87[60] <= result_col87[59];
   result_col87[61] <= result_col87[60];
   result_col87[62] <= result_col87[61];
   result_col87[63] <= result_col87[62];
   result_col87[64] <= result_col87[63];
   result_col87[65] <= result_col87[64];
   result_col87[66] <= result_col87[65];
   result_col87[67] <= result_col87[66];
   result_col87[68] <= result_col87[67];
   result_col87[69] <= result_col87[68];
   result_col87[70] <= result_col87[69];
   result_col87[71] <= result_col87[70];
   result_col87[72] <= result_col87[71];
   result_col87[73] <= result_col87[72];
   result_col87[74] <= result_col87[73];
   result_col87[75] <= result_col87[74];
   result_col87[76] <= result_col87[75];
   result_col87[77] <= result_col87[76];
   result_col87[78] <= result_col87[77];
   result_col87[79] <= result_col87[78];

   result_col88[1] <= data_out_4_88;
   result_col88[2] <= result_col88[1];
   result_col88[3] <= result_col88[2];
   result_col88[4] <= result_col88[3];
   result_col88[5] <= result_col88[4];
   result_col88[6] <= result_col88[5];
   result_col88[7] <= result_col88[6];
   result_col88[8] <= result_col88[7];
   result_col88[9] <= result_col88[8];
   result_col88[10] <= result_col88[9];
   result_col88[11] <= result_col88[10];
   result_col88[12] <= result_col88[11];
   result_col88[13] <= result_col88[12];
   result_col88[14] <= result_col88[13];
   result_col88[15] <= result_col88[14];
   result_col88[16] <= result_col88[15];
   result_col88[17] <= result_col88[16];
   result_col88[18] <= result_col88[17];
   result_col88[19] <= result_col88[18];
   result_col88[20] <= result_col88[19];
   result_col88[21] <= result_col88[20];
   result_col88[22] <= result_col88[21];
   result_col88[23] <= result_col88[22];
   result_col88[24] <= result_col88[23];
   result_col88[25] <= result_col88[24];
   result_col88[26] <= result_col88[25];
   result_col88[27] <= result_col88[26];
   result_col88[28] <= result_col88[27];
   result_col88[29] <= result_col88[28];
   result_col88[30] <= result_col88[29];
   result_col88[31] <= result_col88[30];
   result_col88[32] <= result_col88[31];
   result_col88[33] <= result_col88[32];
   result_col88[34] <= result_col88[33];
   result_col88[35] <= result_col88[34];
   result_col88[36] <= result_col88[35];
   result_col88[37] <= result_col88[36];
   result_col88[38] <= result_col88[37];
   result_col88[39] <= result_col88[38];
   result_col88[40] <= result_col88[39];
   result_col88[41] <= result_col88[40];
   result_col88[42] <= result_col88[41];
   result_col88[43] <= result_col88[42];
   result_col88[44] <= result_col88[43];
   result_col88[45] <= result_col88[44];
   result_col88[46] <= result_col88[45];
   result_col88[47] <= result_col88[46];
   result_col88[48] <= result_col88[47];
   result_col88[49] <= result_col88[48];
   result_col88[50] <= result_col88[49];
   result_col88[51] <= result_col88[50];
   result_col88[52] <= result_col88[51];
   result_col88[53] <= result_col88[52];
   result_col88[54] <= result_col88[53];
   result_col88[55] <= result_col88[54];
   result_col88[56] <= result_col88[55];
   result_col88[57] <= result_col88[56];
   result_col88[58] <= result_col88[57];
   result_col88[59] <= result_col88[58];
   result_col88[60] <= result_col88[59];
   result_col88[61] <= result_col88[60];
   result_col88[62] <= result_col88[61];
   result_col88[63] <= result_col88[62];
   result_col88[64] <= result_col88[63];
   result_col88[65] <= result_col88[64];
   result_col88[66] <= result_col88[65];
   result_col88[67] <= result_col88[66];
   result_col88[68] <= result_col88[67];
   result_col88[69] <= result_col88[68];
   result_col88[70] <= result_col88[69];
   result_col88[71] <= result_col88[70];
   result_col88[72] <= result_col88[71];
   result_col88[73] <= result_col88[72];
   result_col88[74] <= result_col88[73];
   result_col88[75] <= result_col88[74];
   result_col88[76] <= result_col88[75];
   result_col88[77] <= result_col88[76];
   result_col88[78] <= result_col88[77];

   result_col89[1] <= data_out_4_89;
   result_col89[2] <= result_col89[1];
   result_col89[3] <= result_col89[2];
   result_col89[4] <= result_col89[3];
   result_col89[5] <= result_col89[4];
   result_col89[6] <= result_col89[5];
   result_col89[7] <= result_col89[6];
   result_col89[8] <= result_col89[7];
   result_col89[9] <= result_col89[8];
   result_col89[10] <= result_col89[9];
   result_col89[11] <= result_col89[10];
   result_col89[12] <= result_col89[11];
   result_col89[13] <= result_col89[12];
   result_col89[14] <= result_col89[13];
   result_col89[15] <= result_col89[14];
   result_col89[16] <= result_col89[15];
   result_col89[17] <= result_col89[16];
   result_col89[18] <= result_col89[17];
   result_col89[19] <= result_col89[18];
   result_col89[20] <= result_col89[19];
   result_col89[21] <= result_col89[20];
   result_col89[22] <= result_col89[21];
   result_col89[23] <= result_col89[22];
   result_col89[24] <= result_col89[23];
   result_col89[25] <= result_col89[24];
   result_col89[26] <= result_col89[25];
   result_col89[27] <= result_col89[26];
   result_col89[28] <= result_col89[27];
   result_col89[29] <= result_col89[28];
   result_col89[30] <= result_col89[29];
   result_col89[31] <= result_col89[30];
   result_col89[32] <= result_col89[31];
   result_col89[33] <= result_col89[32];
   result_col89[34] <= result_col89[33];
   result_col89[35] <= result_col89[34];
   result_col89[36] <= result_col89[35];
   result_col89[37] <= result_col89[36];
   result_col89[38] <= result_col89[37];
   result_col89[39] <= result_col89[38];
   result_col89[40] <= result_col89[39];
   result_col89[41] <= result_col89[40];
   result_col89[42] <= result_col89[41];
   result_col89[43] <= result_col89[42];
   result_col89[44] <= result_col89[43];
   result_col89[45] <= result_col89[44];
   result_col89[46] <= result_col89[45];
   result_col89[47] <= result_col89[46];
   result_col89[48] <= result_col89[47];
   result_col89[49] <= result_col89[48];
   result_col89[50] <= result_col89[49];
   result_col89[51] <= result_col89[50];
   result_col89[52] <= result_col89[51];
   result_col89[53] <= result_col89[52];
   result_col89[54] <= result_col89[53];
   result_col89[55] <= result_col89[54];
   result_col89[56] <= result_col89[55];
   result_col89[57] <= result_col89[56];
   result_col89[58] <= result_col89[57];
   result_col89[59] <= result_col89[58];
   result_col89[60] <= result_col89[59];
   result_col89[61] <= result_col89[60];
   result_col89[62] <= result_col89[61];
   result_col89[63] <= result_col89[62];
   result_col89[64] <= result_col89[63];
   result_col89[65] <= result_col89[64];
   result_col89[66] <= result_col89[65];
   result_col89[67] <= result_col89[66];
   result_col89[68] <= result_col89[67];
   result_col89[69] <= result_col89[68];
   result_col89[70] <= result_col89[69];
   result_col89[71] <= result_col89[70];
   result_col89[72] <= result_col89[71];
   result_col89[73] <= result_col89[72];
   result_col89[74] <= result_col89[73];
   result_col89[75] <= result_col89[74];
   result_col89[76] <= result_col89[75];
   result_col89[77] <= result_col89[76];

   result_col90[1] <= data_out_4_90;
   result_col90[2] <= result_col90[1];
   result_col90[3] <= result_col90[2];
   result_col90[4] <= result_col90[3];
   result_col90[5] <= result_col90[4];
   result_col90[6] <= result_col90[5];
   result_col90[7] <= result_col90[6];
   result_col90[8] <= result_col90[7];
   result_col90[9] <= result_col90[8];
   result_col90[10] <= result_col90[9];
   result_col90[11] <= result_col90[10];
   result_col90[12] <= result_col90[11];
   result_col90[13] <= result_col90[12];
   result_col90[14] <= result_col90[13];
   result_col90[15] <= result_col90[14];
   result_col90[16] <= result_col90[15];
   result_col90[17] <= result_col90[16];
   result_col90[18] <= result_col90[17];
   result_col90[19] <= result_col90[18];
   result_col90[20] <= result_col90[19];
   result_col90[21] <= result_col90[20];
   result_col90[22] <= result_col90[21];
   result_col90[23] <= result_col90[22];
   result_col90[24] <= result_col90[23];
   result_col90[25] <= result_col90[24];
   result_col90[26] <= result_col90[25];
   result_col90[27] <= result_col90[26];
   result_col90[28] <= result_col90[27];
   result_col90[29] <= result_col90[28];
   result_col90[30] <= result_col90[29];
   result_col90[31] <= result_col90[30];
   result_col90[32] <= result_col90[31];
   result_col90[33] <= result_col90[32];
   result_col90[34] <= result_col90[33];
   result_col90[35] <= result_col90[34];
   result_col90[36] <= result_col90[35];
   result_col90[37] <= result_col90[36];
   result_col90[38] <= result_col90[37];
   result_col90[39] <= result_col90[38];
   result_col90[40] <= result_col90[39];
   result_col90[41] <= result_col90[40];
   result_col90[42] <= result_col90[41];
   result_col90[43] <= result_col90[42];
   result_col90[44] <= result_col90[43];
   result_col90[45] <= result_col90[44];
   result_col90[46] <= result_col90[45];
   result_col90[47] <= result_col90[46];
   result_col90[48] <= result_col90[47];
   result_col90[49] <= result_col90[48];
   result_col90[50] <= result_col90[49];
   result_col90[51] <= result_col90[50];
   result_col90[52] <= result_col90[51];
   result_col90[53] <= result_col90[52];
   result_col90[54] <= result_col90[53];
   result_col90[55] <= result_col90[54];
   result_col90[56] <= result_col90[55];
   result_col90[57] <= result_col90[56];
   result_col90[58] <= result_col90[57];
   result_col90[59] <= result_col90[58];
   result_col90[60] <= result_col90[59];
   result_col90[61] <= result_col90[60];
   result_col90[62] <= result_col90[61];
   result_col90[63] <= result_col90[62];
   result_col90[64] <= result_col90[63];
   result_col90[65] <= result_col90[64];
   result_col90[66] <= result_col90[65];
   result_col90[67] <= result_col90[66];
   result_col90[68] <= result_col90[67];
   result_col90[69] <= result_col90[68];
   result_col90[70] <= result_col90[69];
   result_col90[71] <= result_col90[70];
   result_col90[72] <= result_col90[71];
   result_col90[73] <= result_col90[72];
   result_col90[74] <= result_col90[73];
   result_col90[75] <= result_col90[74];
   result_col90[76] <= result_col90[75];

   result_col91[1] <= data_out_4_91;
   result_col91[2] <= result_col91[1];
   result_col91[3] <= result_col91[2];
   result_col91[4] <= result_col91[3];
   result_col91[5] <= result_col91[4];
   result_col91[6] <= result_col91[5];
   result_col91[7] <= result_col91[6];
   result_col91[8] <= result_col91[7];
   result_col91[9] <= result_col91[8];
   result_col91[10] <= result_col91[9];
   result_col91[11] <= result_col91[10];
   result_col91[12] <= result_col91[11];
   result_col91[13] <= result_col91[12];
   result_col91[14] <= result_col91[13];
   result_col91[15] <= result_col91[14];
   result_col91[16] <= result_col91[15];
   result_col91[17] <= result_col91[16];
   result_col91[18] <= result_col91[17];
   result_col91[19] <= result_col91[18];
   result_col91[20] <= result_col91[19];
   result_col91[21] <= result_col91[20];
   result_col91[22] <= result_col91[21];
   result_col91[23] <= result_col91[22];
   result_col91[24] <= result_col91[23];
   result_col91[25] <= result_col91[24];
   result_col91[26] <= result_col91[25];
   result_col91[27] <= result_col91[26];
   result_col91[28] <= result_col91[27];
   result_col91[29] <= result_col91[28];
   result_col91[30] <= result_col91[29];
   result_col91[31] <= result_col91[30];
   result_col91[32] <= result_col91[31];
   result_col91[33] <= result_col91[32];
   result_col91[34] <= result_col91[33];
   result_col91[35] <= result_col91[34];
   result_col91[36] <= result_col91[35];
   result_col91[37] <= result_col91[36];
   result_col91[38] <= result_col91[37];
   result_col91[39] <= result_col91[38];
   result_col91[40] <= result_col91[39];
   result_col91[41] <= result_col91[40];
   result_col91[42] <= result_col91[41];
   result_col91[43] <= result_col91[42];
   result_col91[44] <= result_col91[43];
   result_col91[45] <= result_col91[44];
   result_col91[46] <= result_col91[45];
   result_col91[47] <= result_col91[46];
   result_col91[48] <= result_col91[47];
   result_col91[49] <= result_col91[48];
   result_col91[50] <= result_col91[49];
   result_col91[51] <= result_col91[50];
   result_col91[52] <= result_col91[51];
   result_col91[53] <= result_col91[52];
   result_col91[54] <= result_col91[53];
   result_col91[55] <= result_col91[54];
   result_col91[56] <= result_col91[55];
   result_col91[57] <= result_col91[56];
   result_col91[58] <= result_col91[57];
   result_col91[59] <= result_col91[58];
   result_col91[60] <= result_col91[59];
   result_col91[61] <= result_col91[60];
   result_col91[62] <= result_col91[61];
   result_col91[63] <= result_col91[62];
   result_col91[64] <= result_col91[63];
   result_col91[65] <= result_col91[64];
   result_col91[66] <= result_col91[65];
   result_col91[67] <= result_col91[66];
   result_col91[68] <= result_col91[67];
   result_col91[69] <= result_col91[68];
   result_col91[70] <= result_col91[69];
   result_col91[71] <= result_col91[70];
   result_col91[72] <= result_col91[71];
   result_col91[73] <= result_col91[72];
   result_col91[74] <= result_col91[73];
   result_col91[75] <= result_col91[74];

   result_col92[1] <= data_out_4_92;
   result_col92[2] <= result_col92[1];
   result_col92[3] <= result_col92[2];
   result_col92[4] <= result_col92[3];
   result_col92[5] <= result_col92[4];
   result_col92[6] <= result_col92[5];
   result_col92[7] <= result_col92[6];
   result_col92[8] <= result_col92[7];
   result_col92[9] <= result_col92[8];
   result_col92[10] <= result_col92[9];
   result_col92[11] <= result_col92[10];
   result_col92[12] <= result_col92[11];
   result_col92[13] <= result_col92[12];
   result_col92[14] <= result_col92[13];
   result_col92[15] <= result_col92[14];
   result_col92[16] <= result_col92[15];
   result_col92[17] <= result_col92[16];
   result_col92[18] <= result_col92[17];
   result_col92[19] <= result_col92[18];
   result_col92[20] <= result_col92[19];
   result_col92[21] <= result_col92[20];
   result_col92[22] <= result_col92[21];
   result_col92[23] <= result_col92[22];
   result_col92[24] <= result_col92[23];
   result_col92[25] <= result_col92[24];
   result_col92[26] <= result_col92[25];
   result_col92[27] <= result_col92[26];
   result_col92[28] <= result_col92[27];
   result_col92[29] <= result_col92[28];
   result_col92[30] <= result_col92[29];
   result_col92[31] <= result_col92[30];
   result_col92[32] <= result_col92[31];
   result_col92[33] <= result_col92[32];
   result_col92[34] <= result_col92[33];
   result_col92[35] <= result_col92[34];
   result_col92[36] <= result_col92[35];
   result_col92[37] <= result_col92[36];
   result_col92[38] <= result_col92[37];
   result_col92[39] <= result_col92[38];
   result_col92[40] <= result_col92[39];
   result_col92[41] <= result_col92[40];
   result_col92[42] <= result_col92[41];
   result_col92[43] <= result_col92[42];
   result_col92[44] <= result_col92[43];
   result_col92[45] <= result_col92[44];
   result_col92[46] <= result_col92[45];
   result_col92[47] <= result_col92[46];
   result_col92[48] <= result_col92[47];
   result_col92[49] <= result_col92[48];
   result_col92[50] <= result_col92[49];
   result_col92[51] <= result_col92[50];
   result_col92[52] <= result_col92[51];
   result_col92[53] <= result_col92[52];
   result_col92[54] <= result_col92[53];
   result_col92[55] <= result_col92[54];
   result_col92[56] <= result_col92[55];
   result_col92[57] <= result_col92[56];
   result_col92[58] <= result_col92[57];
   result_col92[59] <= result_col92[58];
   result_col92[60] <= result_col92[59];
   result_col92[61] <= result_col92[60];
   result_col92[62] <= result_col92[61];
   result_col92[63] <= result_col92[62];
   result_col92[64] <= result_col92[63];
   result_col92[65] <= result_col92[64];
   result_col92[66] <= result_col92[65];
   result_col92[67] <= result_col92[66];
   result_col92[68] <= result_col92[67];
   result_col92[69] <= result_col92[68];
   result_col92[70] <= result_col92[69];
   result_col92[71] <= result_col92[70];
   result_col92[72] <= result_col92[71];
   result_col92[73] <= result_col92[72];
   result_col92[74] <= result_col92[73];

   result_col93[1] <= data_out_4_93;
   result_col93[2] <= result_col93[1];
   result_col93[3] <= result_col93[2];
   result_col93[4] <= result_col93[3];
   result_col93[5] <= result_col93[4];
   result_col93[6] <= result_col93[5];
   result_col93[7] <= result_col93[6];
   result_col93[8] <= result_col93[7];
   result_col93[9] <= result_col93[8];
   result_col93[10] <= result_col93[9];
   result_col93[11] <= result_col93[10];
   result_col93[12] <= result_col93[11];
   result_col93[13] <= result_col93[12];
   result_col93[14] <= result_col93[13];
   result_col93[15] <= result_col93[14];
   result_col93[16] <= result_col93[15];
   result_col93[17] <= result_col93[16];
   result_col93[18] <= result_col93[17];
   result_col93[19] <= result_col93[18];
   result_col93[20] <= result_col93[19];
   result_col93[21] <= result_col93[20];
   result_col93[22] <= result_col93[21];
   result_col93[23] <= result_col93[22];
   result_col93[24] <= result_col93[23];
   result_col93[25] <= result_col93[24];
   result_col93[26] <= result_col93[25];
   result_col93[27] <= result_col93[26];
   result_col93[28] <= result_col93[27];
   result_col93[29] <= result_col93[28];
   result_col93[30] <= result_col93[29];
   result_col93[31] <= result_col93[30];
   result_col93[32] <= result_col93[31];
   result_col93[33] <= result_col93[32];
   result_col93[34] <= result_col93[33];
   result_col93[35] <= result_col93[34];
   result_col93[36] <= result_col93[35];
   result_col93[37] <= result_col93[36];
   result_col93[38] <= result_col93[37];
   result_col93[39] <= result_col93[38];
   result_col93[40] <= result_col93[39];
   result_col93[41] <= result_col93[40];
   result_col93[42] <= result_col93[41];
   result_col93[43] <= result_col93[42];
   result_col93[44] <= result_col93[43];
   result_col93[45] <= result_col93[44];
   result_col93[46] <= result_col93[45];
   result_col93[47] <= result_col93[46];
   result_col93[48] <= result_col93[47];
   result_col93[49] <= result_col93[48];
   result_col93[50] <= result_col93[49];
   result_col93[51] <= result_col93[50];
   result_col93[52] <= result_col93[51];
   result_col93[53] <= result_col93[52];
   result_col93[54] <= result_col93[53];
   result_col93[55] <= result_col93[54];
   result_col93[56] <= result_col93[55];
   result_col93[57] <= result_col93[56];
   result_col93[58] <= result_col93[57];
   result_col93[59] <= result_col93[58];
   result_col93[60] <= result_col93[59];
   result_col93[61] <= result_col93[60];
   result_col93[62] <= result_col93[61];
   result_col93[63] <= result_col93[62];
   result_col93[64] <= result_col93[63];
   result_col93[65] <= result_col93[64];
   result_col93[66] <= result_col93[65];
   result_col93[67] <= result_col93[66];
   result_col93[68] <= result_col93[67];
   result_col93[69] <= result_col93[68];
   result_col93[70] <= result_col93[69];
   result_col93[71] <= result_col93[70];
   result_col93[72] <= result_col93[71];
   result_col93[73] <= result_col93[72];

   result_col94[1] <= data_out_4_94;
   result_col94[2] <= result_col94[1];
   result_col94[3] <= result_col94[2];
   result_col94[4] <= result_col94[3];
   result_col94[5] <= result_col94[4];
   result_col94[6] <= result_col94[5];
   result_col94[7] <= result_col94[6];
   result_col94[8] <= result_col94[7];
   result_col94[9] <= result_col94[8];
   result_col94[10] <= result_col94[9];
   result_col94[11] <= result_col94[10];
   result_col94[12] <= result_col94[11];
   result_col94[13] <= result_col94[12];
   result_col94[14] <= result_col94[13];
   result_col94[15] <= result_col94[14];
   result_col94[16] <= result_col94[15];
   result_col94[17] <= result_col94[16];
   result_col94[18] <= result_col94[17];
   result_col94[19] <= result_col94[18];
   result_col94[20] <= result_col94[19];
   result_col94[21] <= result_col94[20];
   result_col94[22] <= result_col94[21];
   result_col94[23] <= result_col94[22];
   result_col94[24] <= result_col94[23];
   result_col94[25] <= result_col94[24];
   result_col94[26] <= result_col94[25];
   result_col94[27] <= result_col94[26];
   result_col94[28] <= result_col94[27];
   result_col94[29] <= result_col94[28];
   result_col94[30] <= result_col94[29];
   result_col94[31] <= result_col94[30];
   result_col94[32] <= result_col94[31];
   result_col94[33] <= result_col94[32];
   result_col94[34] <= result_col94[33];
   result_col94[35] <= result_col94[34];
   result_col94[36] <= result_col94[35];
   result_col94[37] <= result_col94[36];
   result_col94[38] <= result_col94[37];
   result_col94[39] <= result_col94[38];
   result_col94[40] <= result_col94[39];
   result_col94[41] <= result_col94[40];
   result_col94[42] <= result_col94[41];
   result_col94[43] <= result_col94[42];
   result_col94[44] <= result_col94[43];
   result_col94[45] <= result_col94[44];
   result_col94[46] <= result_col94[45];
   result_col94[47] <= result_col94[46];
   result_col94[48] <= result_col94[47];
   result_col94[49] <= result_col94[48];
   result_col94[50] <= result_col94[49];
   result_col94[51] <= result_col94[50];
   result_col94[52] <= result_col94[51];
   result_col94[53] <= result_col94[52];
   result_col94[54] <= result_col94[53];
   result_col94[55] <= result_col94[54];
   result_col94[56] <= result_col94[55];
   result_col94[57] <= result_col94[56];
   result_col94[58] <= result_col94[57];
   result_col94[59] <= result_col94[58];
   result_col94[60] <= result_col94[59];
   result_col94[61] <= result_col94[60];
   result_col94[62] <= result_col94[61];
   result_col94[63] <= result_col94[62];
   result_col94[64] <= result_col94[63];
   result_col94[65] <= result_col94[64];
   result_col94[66] <= result_col94[65];
   result_col94[67] <= result_col94[66];
   result_col94[68] <= result_col94[67];
   result_col94[69] <= result_col94[68];
   result_col94[70] <= result_col94[69];
   result_col94[71] <= result_col94[70];
   result_col94[72] <= result_col94[71];

   result_col95[1] <= data_out_4_95;
   result_col95[2] <= result_col95[1];
   result_col95[3] <= result_col95[2];
   result_col95[4] <= result_col95[3];
   result_col95[5] <= result_col95[4];
   result_col95[6] <= result_col95[5];
   result_col95[7] <= result_col95[6];
   result_col95[8] <= result_col95[7];
   result_col95[9] <= result_col95[8];
   result_col95[10] <= result_col95[9];
   result_col95[11] <= result_col95[10];
   result_col95[12] <= result_col95[11];
   result_col95[13] <= result_col95[12];
   result_col95[14] <= result_col95[13];
   result_col95[15] <= result_col95[14];
   result_col95[16] <= result_col95[15];
   result_col95[17] <= result_col95[16];
   result_col95[18] <= result_col95[17];
   result_col95[19] <= result_col95[18];
   result_col95[20] <= result_col95[19];
   result_col95[21] <= result_col95[20];
   result_col95[22] <= result_col95[21];
   result_col95[23] <= result_col95[22];
   result_col95[24] <= result_col95[23];
   result_col95[25] <= result_col95[24];
   result_col95[26] <= result_col95[25];
   result_col95[27] <= result_col95[26];
   result_col95[28] <= result_col95[27];
   result_col95[29] <= result_col95[28];
   result_col95[30] <= result_col95[29];
   result_col95[31] <= result_col95[30];
   result_col95[32] <= result_col95[31];
   result_col95[33] <= result_col95[32];
   result_col95[34] <= result_col95[33];
   result_col95[35] <= result_col95[34];
   result_col95[36] <= result_col95[35];
   result_col95[37] <= result_col95[36];
   result_col95[38] <= result_col95[37];
   result_col95[39] <= result_col95[38];
   result_col95[40] <= result_col95[39];
   result_col95[41] <= result_col95[40];
   result_col95[42] <= result_col95[41];
   result_col95[43] <= result_col95[42];
   result_col95[44] <= result_col95[43];
   result_col95[45] <= result_col95[44];
   result_col95[46] <= result_col95[45];
   result_col95[47] <= result_col95[46];
   result_col95[48] <= result_col95[47];
   result_col95[49] <= result_col95[48];
   result_col95[50] <= result_col95[49];
   result_col95[51] <= result_col95[50];
   result_col95[52] <= result_col95[51];
   result_col95[53] <= result_col95[52];
   result_col95[54] <= result_col95[53];
   result_col95[55] <= result_col95[54];
   result_col95[56] <= result_col95[55];
   result_col95[57] <= result_col95[56];
   result_col95[58] <= result_col95[57];
   result_col95[59] <= result_col95[58];
   result_col95[60] <= result_col95[59];
   result_col95[61] <= result_col95[60];
   result_col95[62] <= result_col95[61];
   result_col95[63] <= result_col95[62];
   result_col95[64] <= result_col95[63];
   result_col95[65] <= result_col95[64];
   result_col95[66] <= result_col95[65];
   result_col95[67] <= result_col95[66];
   result_col95[68] <= result_col95[67];
   result_col95[69] <= result_col95[68];
   result_col95[70] <= result_col95[69];
   result_col95[71] <= result_col95[70];

   result_col96[1] <= data_out_4_96;
   result_col96[2] <= result_col96[1];
   result_col96[3] <= result_col96[2];
   result_col96[4] <= result_col96[3];
   result_col96[5] <= result_col96[4];
   result_col96[6] <= result_col96[5];
   result_col96[7] <= result_col96[6];
   result_col96[8] <= result_col96[7];
   result_col96[9] <= result_col96[8];
   result_col96[10] <= result_col96[9];
   result_col96[11] <= result_col96[10];
   result_col96[12] <= result_col96[11];
   result_col96[13] <= result_col96[12];
   result_col96[14] <= result_col96[13];
   result_col96[15] <= result_col96[14];
   result_col96[16] <= result_col96[15];
   result_col96[17] <= result_col96[16];
   result_col96[18] <= result_col96[17];
   result_col96[19] <= result_col96[18];
   result_col96[20] <= result_col96[19];
   result_col96[21] <= result_col96[20];
   result_col96[22] <= result_col96[21];
   result_col96[23] <= result_col96[22];
   result_col96[24] <= result_col96[23];
   result_col96[25] <= result_col96[24];
   result_col96[26] <= result_col96[25];
   result_col96[27] <= result_col96[26];
   result_col96[28] <= result_col96[27];
   result_col96[29] <= result_col96[28];
   result_col96[30] <= result_col96[29];
   result_col96[31] <= result_col96[30];
   result_col96[32] <= result_col96[31];
   result_col96[33] <= result_col96[32];
   result_col96[34] <= result_col96[33];
   result_col96[35] <= result_col96[34];
   result_col96[36] <= result_col96[35];
   result_col96[37] <= result_col96[36];
   result_col96[38] <= result_col96[37];
   result_col96[39] <= result_col96[38];
   result_col96[40] <= result_col96[39];
   result_col96[41] <= result_col96[40];
   result_col96[42] <= result_col96[41];
   result_col96[43] <= result_col96[42];
   result_col96[44] <= result_col96[43];
   result_col96[45] <= result_col96[44];
   result_col96[46] <= result_col96[45];
   result_col96[47] <= result_col96[46];
   result_col96[48] <= result_col96[47];
   result_col96[49] <= result_col96[48];
   result_col96[50] <= result_col96[49];
   result_col96[51] <= result_col96[50];
   result_col96[52] <= result_col96[51];
   result_col96[53] <= result_col96[52];
   result_col96[54] <= result_col96[53];
   result_col96[55] <= result_col96[54];
   result_col96[56] <= result_col96[55];
   result_col96[57] <= result_col96[56];
   result_col96[58] <= result_col96[57];
   result_col96[59] <= result_col96[58];
   result_col96[60] <= result_col96[59];
   result_col96[61] <= result_col96[60];
   result_col96[62] <= result_col96[61];
   result_col96[63] <= result_col96[62];
   result_col96[64] <= result_col96[63];
   result_col96[65] <= result_col96[64];
   result_col96[66] <= result_col96[65];
   result_col96[67] <= result_col96[66];
   result_col96[68] <= result_col96[67];
   result_col96[69] <= result_col96[68];
   result_col96[70] <= result_col96[69];

   result_col97[1] <= data_out_4_97;
   result_col97[2] <= result_col97[1];
   result_col97[3] <= result_col97[2];
   result_col97[4] <= result_col97[3];
   result_col97[5] <= result_col97[4];
   result_col97[6] <= result_col97[5];
   result_col97[7] <= result_col97[6];
   result_col97[8] <= result_col97[7];
   result_col97[9] <= result_col97[8];
   result_col97[10] <= result_col97[9];
   result_col97[11] <= result_col97[10];
   result_col97[12] <= result_col97[11];
   result_col97[13] <= result_col97[12];
   result_col97[14] <= result_col97[13];
   result_col97[15] <= result_col97[14];
   result_col97[16] <= result_col97[15];
   result_col97[17] <= result_col97[16];
   result_col97[18] <= result_col97[17];
   result_col97[19] <= result_col97[18];
   result_col97[20] <= result_col97[19];
   result_col97[21] <= result_col97[20];
   result_col97[22] <= result_col97[21];
   result_col97[23] <= result_col97[22];
   result_col97[24] <= result_col97[23];
   result_col97[25] <= result_col97[24];
   result_col97[26] <= result_col97[25];
   result_col97[27] <= result_col97[26];
   result_col97[28] <= result_col97[27];
   result_col97[29] <= result_col97[28];
   result_col97[30] <= result_col97[29];
   result_col97[31] <= result_col97[30];
   result_col97[32] <= result_col97[31];
   result_col97[33] <= result_col97[32];
   result_col97[34] <= result_col97[33];
   result_col97[35] <= result_col97[34];
   result_col97[36] <= result_col97[35];
   result_col97[37] <= result_col97[36];
   result_col97[38] <= result_col97[37];
   result_col97[39] <= result_col97[38];
   result_col97[40] <= result_col97[39];
   result_col97[41] <= result_col97[40];
   result_col97[42] <= result_col97[41];
   result_col97[43] <= result_col97[42];
   result_col97[44] <= result_col97[43];
   result_col97[45] <= result_col97[44];
   result_col97[46] <= result_col97[45];
   result_col97[47] <= result_col97[46];
   result_col97[48] <= result_col97[47];
   result_col97[49] <= result_col97[48];
   result_col97[50] <= result_col97[49];
   result_col97[51] <= result_col97[50];
   result_col97[52] <= result_col97[51];
   result_col97[53] <= result_col97[52];
   result_col97[54] <= result_col97[53];
   result_col97[55] <= result_col97[54];
   result_col97[56] <= result_col97[55];
   result_col97[57] <= result_col97[56];
   result_col97[58] <= result_col97[57];
   result_col97[59] <= result_col97[58];
   result_col97[60] <= result_col97[59];
   result_col97[61] <= result_col97[60];
   result_col97[62] <= result_col97[61];
   result_col97[63] <= result_col97[62];
   result_col97[64] <= result_col97[63];
   result_col97[65] <= result_col97[64];
   result_col97[66] <= result_col97[65];
   result_col97[67] <= result_col97[66];
   result_col97[68] <= result_col97[67];
   result_col97[69] <= result_col97[68];

   result_col98[1] <= data_out_4_98;
   result_col98[2] <= result_col98[1];
   result_col98[3] <= result_col98[2];
   result_col98[4] <= result_col98[3];
   result_col98[5] <= result_col98[4];
   result_col98[6] <= result_col98[5];
   result_col98[7] <= result_col98[6];
   result_col98[8] <= result_col98[7];
   result_col98[9] <= result_col98[8];
   result_col98[10] <= result_col98[9];
   result_col98[11] <= result_col98[10];
   result_col98[12] <= result_col98[11];
   result_col98[13] <= result_col98[12];
   result_col98[14] <= result_col98[13];
   result_col98[15] <= result_col98[14];
   result_col98[16] <= result_col98[15];
   result_col98[17] <= result_col98[16];
   result_col98[18] <= result_col98[17];
   result_col98[19] <= result_col98[18];
   result_col98[20] <= result_col98[19];
   result_col98[21] <= result_col98[20];
   result_col98[22] <= result_col98[21];
   result_col98[23] <= result_col98[22];
   result_col98[24] <= result_col98[23];
   result_col98[25] <= result_col98[24];
   result_col98[26] <= result_col98[25];
   result_col98[27] <= result_col98[26];
   result_col98[28] <= result_col98[27];
   result_col98[29] <= result_col98[28];
   result_col98[30] <= result_col98[29];
   result_col98[31] <= result_col98[30];
   result_col98[32] <= result_col98[31];
   result_col98[33] <= result_col98[32];
   result_col98[34] <= result_col98[33];
   result_col98[35] <= result_col98[34];
   result_col98[36] <= result_col98[35];
   result_col98[37] <= result_col98[36];
   result_col98[38] <= result_col98[37];
   result_col98[39] <= result_col98[38];
   result_col98[40] <= result_col98[39];
   result_col98[41] <= result_col98[40];
   result_col98[42] <= result_col98[41];
   result_col98[43] <= result_col98[42];
   result_col98[44] <= result_col98[43];
   result_col98[45] <= result_col98[44];
   result_col98[46] <= result_col98[45];
   result_col98[47] <= result_col98[46];
   result_col98[48] <= result_col98[47];
   result_col98[49] <= result_col98[48];
   result_col98[50] <= result_col98[49];
   result_col98[51] <= result_col98[50];
   result_col98[52] <= result_col98[51];
   result_col98[53] <= result_col98[52];
   result_col98[54] <= result_col98[53];
   result_col98[55] <= result_col98[54];
   result_col98[56] <= result_col98[55];
   result_col98[57] <= result_col98[56];
   result_col98[58] <= result_col98[57];
   result_col98[59] <= result_col98[58];
   result_col98[60] <= result_col98[59];
   result_col98[61] <= result_col98[60];
   result_col98[62] <= result_col98[61];
   result_col98[63] <= result_col98[62];
   result_col98[64] <= result_col98[63];
   result_col98[65] <= result_col98[64];
   result_col98[66] <= result_col98[65];
   result_col98[67] <= result_col98[66];
   result_col98[68] <= result_col98[67];

   result_col99[1] <= data_out_4_99;
   result_col99[2] <= result_col99[1];
   result_col99[3] <= result_col99[2];
   result_col99[4] <= result_col99[3];
   result_col99[5] <= result_col99[4];
   result_col99[6] <= result_col99[5];
   result_col99[7] <= result_col99[6];
   result_col99[8] <= result_col99[7];
   result_col99[9] <= result_col99[8];
   result_col99[10] <= result_col99[9];
   result_col99[11] <= result_col99[10];
   result_col99[12] <= result_col99[11];
   result_col99[13] <= result_col99[12];
   result_col99[14] <= result_col99[13];
   result_col99[15] <= result_col99[14];
   result_col99[16] <= result_col99[15];
   result_col99[17] <= result_col99[16];
   result_col99[18] <= result_col99[17];
   result_col99[19] <= result_col99[18];
   result_col99[20] <= result_col99[19];
   result_col99[21] <= result_col99[20];
   result_col99[22] <= result_col99[21];
   result_col99[23] <= result_col99[22];
   result_col99[24] <= result_col99[23];
   result_col99[25] <= result_col99[24];
   result_col99[26] <= result_col99[25];
   result_col99[27] <= result_col99[26];
   result_col99[28] <= result_col99[27];
   result_col99[29] <= result_col99[28];
   result_col99[30] <= result_col99[29];
   result_col99[31] <= result_col99[30];
   result_col99[32] <= result_col99[31];
   result_col99[33] <= result_col99[32];
   result_col99[34] <= result_col99[33];
   result_col99[35] <= result_col99[34];
   result_col99[36] <= result_col99[35];
   result_col99[37] <= result_col99[36];
   result_col99[38] <= result_col99[37];
   result_col99[39] <= result_col99[38];
   result_col99[40] <= result_col99[39];
   result_col99[41] <= result_col99[40];
   result_col99[42] <= result_col99[41];
   result_col99[43] <= result_col99[42];
   result_col99[44] <= result_col99[43];
   result_col99[45] <= result_col99[44];
   result_col99[46] <= result_col99[45];
   result_col99[47] <= result_col99[46];
   result_col99[48] <= result_col99[47];
   result_col99[49] <= result_col99[48];
   result_col99[50] <= result_col99[49];
   result_col99[51] <= result_col99[50];
   result_col99[52] <= result_col99[51];
   result_col99[53] <= result_col99[52];
   result_col99[54] <= result_col99[53];
   result_col99[55] <= result_col99[54];
   result_col99[56] <= result_col99[55];
   result_col99[57] <= result_col99[56];
   result_col99[58] <= result_col99[57];
   result_col99[59] <= result_col99[58];
   result_col99[60] <= result_col99[59];
   result_col99[61] <= result_col99[60];
   result_col99[62] <= result_col99[61];
   result_col99[63] <= result_col99[62];
   result_col99[64] <= result_col99[63];
   result_col99[65] <= result_col99[64];
   result_col99[66] <= result_col99[65];
   result_col99[67] <= result_col99[66];

   result_col100[1] <= data_out_4_100;
   result_col100[2] <= result_col100[1];
   result_col100[3] <= result_col100[2];
   result_col100[4] <= result_col100[3];
   result_col100[5] <= result_col100[4];
   result_col100[6] <= result_col100[5];
   result_col100[7] <= result_col100[6];
   result_col100[8] <= result_col100[7];
   result_col100[9] <= result_col100[8];
   result_col100[10] <= result_col100[9];
   result_col100[11] <= result_col100[10];
   result_col100[12] <= result_col100[11];
   result_col100[13] <= result_col100[12];
   result_col100[14] <= result_col100[13];
   result_col100[15] <= result_col100[14];
   result_col100[16] <= result_col100[15];
   result_col100[17] <= result_col100[16];
   result_col100[18] <= result_col100[17];
   result_col100[19] <= result_col100[18];
   result_col100[20] <= result_col100[19];
   result_col100[21] <= result_col100[20];
   result_col100[22] <= result_col100[21];
   result_col100[23] <= result_col100[22];
   result_col100[24] <= result_col100[23];
   result_col100[25] <= result_col100[24];
   result_col100[26] <= result_col100[25];
   result_col100[27] <= result_col100[26];
   result_col100[28] <= result_col100[27];
   result_col100[29] <= result_col100[28];
   result_col100[30] <= result_col100[29];
   result_col100[31] <= result_col100[30];
   result_col100[32] <= result_col100[31];
   result_col100[33] <= result_col100[32];
   result_col100[34] <= result_col100[33];
   result_col100[35] <= result_col100[34];
   result_col100[36] <= result_col100[35];
   result_col100[37] <= result_col100[36];
   result_col100[38] <= result_col100[37];
   result_col100[39] <= result_col100[38];
   result_col100[40] <= result_col100[39];
   result_col100[41] <= result_col100[40];
   result_col100[42] <= result_col100[41];
   result_col100[43] <= result_col100[42];
   result_col100[44] <= result_col100[43];
   result_col100[45] <= result_col100[44];
   result_col100[46] <= result_col100[45];
   result_col100[47] <= result_col100[46];
   result_col100[48] <= result_col100[47];
   result_col100[49] <= result_col100[48];
   result_col100[50] <= result_col100[49];
   result_col100[51] <= result_col100[50];
   result_col100[52] <= result_col100[51];
   result_col100[53] <= result_col100[52];
   result_col100[54] <= result_col100[53];
   result_col100[55] <= result_col100[54];
   result_col100[56] <= result_col100[55];
   result_col100[57] <= result_col100[56];
   result_col100[58] <= result_col100[57];
   result_col100[59] <= result_col100[58];
   result_col100[60] <= result_col100[59];
   result_col100[61] <= result_col100[60];
   result_col100[62] <= result_col100[61];
   result_col100[63] <= result_col100[62];
   result_col100[64] <= result_col100[63];
   result_col100[65] <= result_col100[64];
   result_col100[66] <= result_col100[65];

   result_col101[1] <= data_out_4_101;
   result_col101[2] <= result_col101[1];
   result_col101[3] <= result_col101[2];
   result_col101[4] <= result_col101[3];
   result_col101[5] <= result_col101[4];
   result_col101[6] <= result_col101[5];
   result_col101[7] <= result_col101[6];
   result_col101[8] <= result_col101[7];
   result_col101[9] <= result_col101[8];
   result_col101[10] <= result_col101[9];
   result_col101[11] <= result_col101[10];
   result_col101[12] <= result_col101[11];
   result_col101[13] <= result_col101[12];
   result_col101[14] <= result_col101[13];
   result_col101[15] <= result_col101[14];
   result_col101[16] <= result_col101[15];
   result_col101[17] <= result_col101[16];
   result_col101[18] <= result_col101[17];
   result_col101[19] <= result_col101[18];
   result_col101[20] <= result_col101[19];
   result_col101[21] <= result_col101[20];
   result_col101[22] <= result_col101[21];
   result_col101[23] <= result_col101[22];
   result_col101[24] <= result_col101[23];
   result_col101[25] <= result_col101[24];
   result_col101[26] <= result_col101[25];
   result_col101[27] <= result_col101[26];
   result_col101[28] <= result_col101[27];
   result_col101[29] <= result_col101[28];
   result_col101[30] <= result_col101[29];
   result_col101[31] <= result_col101[30];
   result_col101[32] <= result_col101[31];
   result_col101[33] <= result_col101[32];
   result_col101[34] <= result_col101[33];
   result_col101[35] <= result_col101[34];
   result_col101[36] <= result_col101[35];
   result_col101[37] <= result_col101[36];
   result_col101[38] <= result_col101[37];
   result_col101[39] <= result_col101[38];
   result_col101[40] <= result_col101[39];
   result_col101[41] <= result_col101[40];
   result_col101[42] <= result_col101[41];
   result_col101[43] <= result_col101[42];
   result_col101[44] <= result_col101[43];
   result_col101[45] <= result_col101[44];
   result_col101[46] <= result_col101[45];
   result_col101[47] <= result_col101[46];
   result_col101[48] <= result_col101[47];
   result_col101[49] <= result_col101[48];
   result_col101[50] <= result_col101[49];
   result_col101[51] <= result_col101[50];
   result_col101[52] <= result_col101[51];
   result_col101[53] <= result_col101[52];
   result_col101[54] <= result_col101[53];
   result_col101[55] <= result_col101[54];
   result_col101[56] <= result_col101[55];
   result_col101[57] <= result_col101[56];
   result_col101[58] <= result_col101[57];
   result_col101[59] <= result_col101[58];
   result_col101[60] <= result_col101[59];
   result_col101[61] <= result_col101[60];
   result_col101[62] <= result_col101[61];
   result_col101[63] <= result_col101[62];
   result_col101[64] <= result_col101[63];
   result_col101[65] <= result_col101[64];

   result_col102[1] <= data_out_4_102;
   result_col102[2] <= result_col102[1];
   result_col102[3] <= result_col102[2];
   result_col102[4] <= result_col102[3];
   result_col102[5] <= result_col102[4];
   result_col102[6] <= result_col102[5];
   result_col102[7] <= result_col102[6];
   result_col102[8] <= result_col102[7];
   result_col102[9] <= result_col102[8];
   result_col102[10] <= result_col102[9];
   result_col102[11] <= result_col102[10];
   result_col102[12] <= result_col102[11];
   result_col102[13] <= result_col102[12];
   result_col102[14] <= result_col102[13];
   result_col102[15] <= result_col102[14];
   result_col102[16] <= result_col102[15];
   result_col102[17] <= result_col102[16];
   result_col102[18] <= result_col102[17];
   result_col102[19] <= result_col102[18];
   result_col102[20] <= result_col102[19];
   result_col102[21] <= result_col102[20];
   result_col102[22] <= result_col102[21];
   result_col102[23] <= result_col102[22];
   result_col102[24] <= result_col102[23];
   result_col102[25] <= result_col102[24];
   result_col102[26] <= result_col102[25];
   result_col102[27] <= result_col102[26];
   result_col102[28] <= result_col102[27];
   result_col102[29] <= result_col102[28];
   result_col102[30] <= result_col102[29];
   result_col102[31] <= result_col102[30];
   result_col102[32] <= result_col102[31];
   result_col102[33] <= result_col102[32];
   result_col102[34] <= result_col102[33];
   result_col102[35] <= result_col102[34];
   result_col102[36] <= result_col102[35];
   result_col102[37] <= result_col102[36];
   result_col102[38] <= result_col102[37];
   result_col102[39] <= result_col102[38];
   result_col102[40] <= result_col102[39];
   result_col102[41] <= result_col102[40];
   result_col102[42] <= result_col102[41];
   result_col102[43] <= result_col102[42];
   result_col102[44] <= result_col102[43];
   result_col102[45] <= result_col102[44];
   result_col102[46] <= result_col102[45];
   result_col102[47] <= result_col102[46];
   result_col102[48] <= result_col102[47];
   result_col102[49] <= result_col102[48];
   result_col102[50] <= result_col102[49];
   result_col102[51] <= result_col102[50];
   result_col102[52] <= result_col102[51];
   result_col102[53] <= result_col102[52];
   result_col102[54] <= result_col102[53];
   result_col102[55] <= result_col102[54];
   result_col102[56] <= result_col102[55];
   result_col102[57] <= result_col102[56];
   result_col102[58] <= result_col102[57];
   result_col102[59] <= result_col102[58];
   result_col102[60] <= result_col102[59];
   result_col102[61] <= result_col102[60];
   result_col102[62] <= result_col102[61];
   result_col102[63] <= result_col102[62];
   result_col102[64] <= result_col102[63];

   result_col103[1] <= data_out_4_103;
   result_col103[2] <= result_col103[1];
   result_col103[3] <= result_col103[2];
   result_col103[4] <= result_col103[3];
   result_col103[5] <= result_col103[4];
   result_col103[6] <= result_col103[5];
   result_col103[7] <= result_col103[6];
   result_col103[8] <= result_col103[7];
   result_col103[9] <= result_col103[8];
   result_col103[10] <= result_col103[9];
   result_col103[11] <= result_col103[10];
   result_col103[12] <= result_col103[11];
   result_col103[13] <= result_col103[12];
   result_col103[14] <= result_col103[13];
   result_col103[15] <= result_col103[14];
   result_col103[16] <= result_col103[15];
   result_col103[17] <= result_col103[16];
   result_col103[18] <= result_col103[17];
   result_col103[19] <= result_col103[18];
   result_col103[20] <= result_col103[19];
   result_col103[21] <= result_col103[20];
   result_col103[22] <= result_col103[21];
   result_col103[23] <= result_col103[22];
   result_col103[24] <= result_col103[23];
   result_col103[25] <= result_col103[24];
   result_col103[26] <= result_col103[25];
   result_col103[27] <= result_col103[26];
   result_col103[28] <= result_col103[27];
   result_col103[29] <= result_col103[28];
   result_col103[30] <= result_col103[29];
   result_col103[31] <= result_col103[30];
   result_col103[32] <= result_col103[31];
   result_col103[33] <= result_col103[32];
   result_col103[34] <= result_col103[33];
   result_col103[35] <= result_col103[34];
   result_col103[36] <= result_col103[35];
   result_col103[37] <= result_col103[36];
   result_col103[38] <= result_col103[37];
   result_col103[39] <= result_col103[38];
   result_col103[40] <= result_col103[39];
   result_col103[41] <= result_col103[40];
   result_col103[42] <= result_col103[41];
   result_col103[43] <= result_col103[42];
   result_col103[44] <= result_col103[43];
   result_col103[45] <= result_col103[44];
   result_col103[46] <= result_col103[45];
   result_col103[47] <= result_col103[46];
   result_col103[48] <= result_col103[47];
   result_col103[49] <= result_col103[48];
   result_col103[50] <= result_col103[49];
   result_col103[51] <= result_col103[50];
   result_col103[52] <= result_col103[51];
   result_col103[53] <= result_col103[52];
   result_col103[54] <= result_col103[53];
   result_col103[55] <= result_col103[54];
   result_col103[56] <= result_col103[55];
   result_col103[57] <= result_col103[56];
   result_col103[58] <= result_col103[57];
   result_col103[59] <= result_col103[58];
   result_col103[60] <= result_col103[59];
   result_col103[61] <= result_col103[60];
   result_col103[62] <= result_col103[61];
   result_col103[63] <= result_col103[62];

   result_col104[1] <= data_out_4_104;
   result_col104[2] <= result_col104[1];
   result_col104[3] <= result_col104[2];
   result_col104[4] <= result_col104[3];
   result_col104[5] <= result_col104[4];
   result_col104[6] <= result_col104[5];
   result_col104[7] <= result_col104[6];
   result_col104[8] <= result_col104[7];
   result_col104[9] <= result_col104[8];
   result_col104[10] <= result_col104[9];
   result_col104[11] <= result_col104[10];
   result_col104[12] <= result_col104[11];
   result_col104[13] <= result_col104[12];
   result_col104[14] <= result_col104[13];
   result_col104[15] <= result_col104[14];
   result_col104[16] <= result_col104[15];
   result_col104[17] <= result_col104[16];
   result_col104[18] <= result_col104[17];
   result_col104[19] <= result_col104[18];
   result_col104[20] <= result_col104[19];
   result_col104[21] <= result_col104[20];
   result_col104[22] <= result_col104[21];
   result_col104[23] <= result_col104[22];
   result_col104[24] <= result_col104[23];
   result_col104[25] <= result_col104[24];
   result_col104[26] <= result_col104[25];
   result_col104[27] <= result_col104[26];
   result_col104[28] <= result_col104[27];
   result_col104[29] <= result_col104[28];
   result_col104[30] <= result_col104[29];
   result_col104[31] <= result_col104[30];
   result_col104[32] <= result_col104[31];
   result_col104[33] <= result_col104[32];
   result_col104[34] <= result_col104[33];
   result_col104[35] <= result_col104[34];
   result_col104[36] <= result_col104[35];
   result_col104[37] <= result_col104[36];
   result_col104[38] <= result_col104[37];
   result_col104[39] <= result_col104[38];
   result_col104[40] <= result_col104[39];
   result_col104[41] <= result_col104[40];
   result_col104[42] <= result_col104[41];
   result_col104[43] <= result_col104[42];
   result_col104[44] <= result_col104[43];
   result_col104[45] <= result_col104[44];
   result_col104[46] <= result_col104[45];
   result_col104[47] <= result_col104[46];
   result_col104[48] <= result_col104[47];
   result_col104[49] <= result_col104[48];
   result_col104[50] <= result_col104[49];
   result_col104[51] <= result_col104[50];
   result_col104[52] <= result_col104[51];
   result_col104[53] <= result_col104[52];
   result_col104[54] <= result_col104[53];
   result_col104[55] <= result_col104[54];
   result_col104[56] <= result_col104[55];
   result_col104[57] <= result_col104[56];
   result_col104[58] <= result_col104[57];
   result_col104[59] <= result_col104[58];
   result_col104[60] <= result_col104[59];
   result_col104[61] <= result_col104[60];
   result_col104[62] <= result_col104[61];

   result_col105[1] <= data_out_4_105;
   result_col105[2] <= result_col105[1];
   result_col105[3] <= result_col105[2];
   result_col105[4] <= result_col105[3];
   result_col105[5] <= result_col105[4];
   result_col105[6] <= result_col105[5];
   result_col105[7] <= result_col105[6];
   result_col105[8] <= result_col105[7];
   result_col105[9] <= result_col105[8];
   result_col105[10] <= result_col105[9];
   result_col105[11] <= result_col105[10];
   result_col105[12] <= result_col105[11];
   result_col105[13] <= result_col105[12];
   result_col105[14] <= result_col105[13];
   result_col105[15] <= result_col105[14];
   result_col105[16] <= result_col105[15];
   result_col105[17] <= result_col105[16];
   result_col105[18] <= result_col105[17];
   result_col105[19] <= result_col105[18];
   result_col105[20] <= result_col105[19];
   result_col105[21] <= result_col105[20];
   result_col105[22] <= result_col105[21];
   result_col105[23] <= result_col105[22];
   result_col105[24] <= result_col105[23];
   result_col105[25] <= result_col105[24];
   result_col105[26] <= result_col105[25];
   result_col105[27] <= result_col105[26];
   result_col105[28] <= result_col105[27];
   result_col105[29] <= result_col105[28];
   result_col105[30] <= result_col105[29];
   result_col105[31] <= result_col105[30];
   result_col105[32] <= result_col105[31];
   result_col105[33] <= result_col105[32];
   result_col105[34] <= result_col105[33];
   result_col105[35] <= result_col105[34];
   result_col105[36] <= result_col105[35];
   result_col105[37] <= result_col105[36];
   result_col105[38] <= result_col105[37];
   result_col105[39] <= result_col105[38];
   result_col105[40] <= result_col105[39];
   result_col105[41] <= result_col105[40];
   result_col105[42] <= result_col105[41];
   result_col105[43] <= result_col105[42];
   result_col105[44] <= result_col105[43];
   result_col105[45] <= result_col105[44];
   result_col105[46] <= result_col105[45];
   result_col105[47] <= result_col105[46];
   result_col105[48] <= result_col105[47];
   result_col105[49] <= result_col105[48];
   result_col105[50] <= result_col105[49];
   result_col105[51] <= result_col105[50];
   result_col105[52] <= result_col105[51];
   result_col105[53] <= result_col105[52];
   result_col105[54] <= result_col105[53];
   result_col105[55] <= result_col105[54];
   result_col105[56] <= result_col105[55];
   result_col105[57] <= result_col105[56];
   result_col105[58] <= result_col105[57];
   result_col105[59] <= result_col105[58];
   result_col105[60] <= result_col105[59];
   result_col105[61] <= result_col105[60];

   result_col106[1] <= data_out_4_106;
   result_col106[2] <= result_col106[1];
   result_col106[3] <= result_col106[2];
   result_col106[4] <= result_col106[3];
   result_col106[5] <= result_col106[4];
   result_col106[6] <= result_col106[5];
   result_col106[7] <= result_col106[6];
   result_col106[8] <= result_col106[7];
   result_col106[9] <= result_col106[8];
   result_col106[10] <= result_col106[9];
   result_col106[11] <= result_col106[10];
   result_col106[12] <= result_col106[11];
   result_col106[13] <= result_col106[12];
   result_col106[14] <= result_col106[13];
   result_col106[15] <= result_col106[14];
   result_col106[16] <= result_col106[15];
   result_col106[17] <= result_col106[16];
   result_col106[18] <= result_col106[17];
   result_col106[19] <= result_col106[18];
   result_col106[20] <= result_col106[19];
   result_col106[21] <= result_col106[20];
   result_col106[22] <= result_col106[21];
   result_col106[23] <= result_col106[22];
   result_col106[24] <= result_col106[23];
   result_col106[25] <= result_col106[24];
   result_col106[26] <= result_col106[25];
   result_col106[27] <= result_col106[26];
   result_col106[28] <= result_col106[27];
   result_col106[29] <= result_col106[28];
   result_col106[30] <= result_col106[29];
   result_col106[31] <= result_col106[30];
   result_col106[32] <= result_col106[31];
   result_col106[33] <= result_col106[32];
   result_col106[34] <= result_col106[33];
   result_col106[35] <= result_col106[34];
   result_col106[36] <= result_col106[35];
   result_col106[37] <= result_col106[36];
   result_col106[38] <= result_col106[37];
   result_col106[39] <= result_col106[38];
   result_col106[40] <= result_col106[39];
   result_col106[41] <= result_col106[40];
   result_col106[42] <= result_col106[41];
   result_col106[43] <= result_col106[42];
   result_col106[44] <= result_col106[43];
   result_col106[45] <= result_col106[44];
   result_col106[46] <= result_col106[45];
   result_col106[47] <= result_col106[46];
   result_col106[48] <= result_col106[47];
   result_col106[49] <= result_col106[48];
   result_col106[50] <= result_col106[49];
   result_col106[51] <= result_col106[50];
   result_col106[52] <= result_col106[51];
   result_col106[53] <= result_col106[52];
   result_col106[54] <= result_col106[53];
   result_col106[55] <= result_col106[54];
   result_col106[56] <= result_col106[55];
   result_col106[57] <= result_col106[56];
   result_col106[58] <= result_col106[57];
   result_col106[59] <= result_col106[58];
   result_col106[60] <= result_col106[59];

   result_col107[1] <= data_out_4_107;
   result_col107[2] <= result_col107[1];
   result_col107[3] <= result_col107[2];
   result_col107[4] <= result_col107[3];
   result_col107[5] <= result_col107[4];
   result_col107[6] <= result_col107[5];
   result_col107[7] <= result_col107[6];
   result_col107[8] <= result_col107[7];
   result_col107[9] <= result_col107[8];
   result_col107[10] <= result_col107[9];
   result_col107[11] <= result_col107[10];
   result_col107[12] <= result_col107[11];
   result_col107[13] <= result_col107[12];
   result_col107[14] <= result_col107[13];
   result_col107[15] <= result_col107[14];
   result_col107[16] <= result_col107[15];
   result_col107[17] <= result_col107[16];
   result_col107[18] <= result_col107[17];
   result_col107[19] <= result_col107[18];
   result_col107[20] <= result_col107[19];
   result_col107[21] <= result_col107[20];
   result_col107[22] <= result_col107[21];
   result_col107[23] <= result_col107[22];
   result_col107[24] <= result_col107[23];
   result_col107[25] <= result_col107[24];
   result_col107[26] <= result_col107[25];
   result_col107[27] <= result_col107[26];
   result_col107[28] <= result_col107[27];
   result_col107[29] <= result_col107[28];
   result_col107[30] <= result_col107[29];
   result_col107[31] <= result_col107[30];
   result_col107[32] <= result_col107[31];
   result_col107[33] <= result_col107[32];
   result_col107[34] <= result_col107[33];
   result_col107[35] <= result_col107[34];
   result_col107[36] <= result_col107[35];
   result_col107[37] <= result_col107[36];
   result_col107[38] <= result_col107[37];
   result_col107[39] <= result_col107[38];
   result_col107[40] <= result_col107[39];
   result_col107[41] <= result_col107[40];
   result_col107[42] <= result_col107[41];
   result_col107[43] <= result_col107[42];
   result_col107[44] <= result_col107[43];
   result_col107[45] <= result_col107[44];
   result_col107[46] <= result_col107[45];
   result_col107[47] <= result_col107[46];
   result_col107[48] <= result_col107[47];
   result_col107[49] <= result_col107[48];
   result_col107[50] <= result_col107[49];
   result_col107[51] <= result_col107[50];
   result_col107[52] <= result_col107[51];
   result_col107[53] <= result_col107[52];
   result_col107[54] <= result_col107[53];
   result_col107[55] <= result_col107[54];
   result_col107[56] <= result_col107[55];
   result_col107[57] <= result_col107[56];
   result_col107[58] <= result_col107[57];
   result_col107[59] <= result_col107[58];

   result_col108[1] <= data_out_4_108;
   result_col108[2] <= result_col108[1];
   result_col108[3] <= result_col108[2];
   result_col108[4] <= result_col108[3];
   result_col108[5] <= result_col108[4];
   result_col108[6] <= result_col108[5];
   result_col108[7] <= result_col108[6];
   result_col108[8] <= result_col108[7];
   result_col108[9] <= result_col108[8];
   result_col108[10] <= result_col108[9];
   result_col108[11] <= result_col108[10];
   result_col108[12] <= result_col108[11];
   result_col108[13] <= result_col108[12];
   result_col108[14] <= result_col108[13];
   result_col108[15] <= result_col108[14];
   result_col108[16] <= result_col108[15];
   result_col108[17] <= result_col108[16];
   result_col108[18] <= result_col108[17];
   result_col108[19] <= result_col108[18];
   result_col108[20] <= result_col108[19];
   result_col108[21] <= result_col108[20];
   result_col108[22] <= result_col108[21];
   result_col108[23] <= result_col108[22];
   result_col108[24] <= result_col108[23];
   result_col108[25] <= result_col108[24];
   result_col108[26] <= result_col108[25];
   result_col108[27] <= result_col108[26];
   result_col108[28] <= result_col108[27];
   result_col108[29] <= result_col108[28];
   result_col108[30] <= result_col108[29];
   result_col108[31] <= result_col108[30];
   result_col108[32] <= result_col108[31];
   result_col108[33] <= result_col108[32];
   result_col108[34] <= result_col108[33];
   result_col108[35] <= result_col108[34];
   result_col108[36] <= result_col108[35];
   result_col108[37] <= result_col108[36];
   result_col108[38] <= result_col108[37];
   result_col108[39] <= result_col108[38];
   result_col108[40] <= result_col108[39];
   result_col108[41] <= result_col108[40];
   result_col108[42] <= result_col108[41];
   result_col108[43] <= result_col108[42];
   result_col108[44] <= result_col108[43];
   result_col108[45] <= result_col108[44];
   result_col108[46] <= result_col108[45];
   result_col108[47] <= result_col108[46];
   result_col108[48] <= result_col108[47];
   result_col108[49] <= result_col108[48];
   result_col108[50] <= result_col108[49];
   result_col108[51] <= result_col108[50];
   result_col108[52] <= result_col108[51];
   result_col108[53] <= result_col108[52];
   result_col108[54] <= result_col108[53];
   result_col108[55] <= result_col108[54];
   result_col108[56] <= result_col108[55];
   result_col108[57] <= result_col108[56];
   result_col108[58] <= result_col108[57];

   result_col109[1] <= data_out_4_109;
   result_col109[2] <= result_col109[1];
   result_col109[3] <= result_col109[2];
   result_col109[4] <= result_col109[3];
   result_col109[5] <= result_col109[4];
   result_col109[6] <= result_col109[5];
   result_col109[7] <= result_col109[6];
   result_col109[8] <= result_col109[7];
   result_col109[9] <= result_col109[8];
   result_col109[10] <= result_col109[9];
   result_col109[11] <= result_col109[10];
   result_col109[12] <= result_col109[11];
   result_col109[13] <= result_col109[12];
   result_col109[14] <= result_col109[13];
   result_col109[15] <= result_col109[14];
   result_col109[16] <= result_col109[15];
   result_col109[17] <= result_col109[16];
   result_col109[18] <= result_col109[17];
   result_col109[19] <= result_col109[18];
   result_col109[20] <= result_col109[19];
   result_col109[21] <= result_col109[20];
   result_col109[22] <= result_col109[21];
   result_col109[23] <= result_col109[22];
   result_col109[24] <= result_col109[23];
   result_col109[25] <= result_col109[24];
   result_col109[26] <= result_col109[25];
   result_col109[27] <= result_col109[26];
   result_col109[28] <= result_col109[27];
   result_col109[29] <= result_col109[28];
   result_col109[30] <= result_col109[29];
   result_col109[31] <= result_col109[30];
   result_col109[32] <= result_col109[31];
   result_col109[33] <= result_col109[32];
   result_col109[34] <= result_col109[33];
   result_col109[35] <= result_col109[34];
   result_col109[36] <= result_col109[35];
   result_col109[37] <= result_col109[36];
   result_col109[38] <= result_col109[37];
   result_col109[39] <= result_col109[38];
   result_col109[40] <= result_col109[39];
   result_col109[41] <= result_col109[40];
   result_col109[42] <= result_col109[41];
   result_col109[43] <= result_col109[42];
   result_col109[44] <= result_col109[43];
   result_col109[45] <= result_col109[44];
   result_col109[46] <= result_col109[45];
   result_col109[47] <= result_col109[46];
   result_col109[48] <= result_col109[47];
   result_col109[49] <= result_col109[48];
   result_col109[50] <= result_col109[49];
   result_col109[51] <= result_col109[50];
   result_col109[52] <= result_col109[51];
   result_col109[53] <= result_col109[52];
   result_col109[54] <= result_col109[53];
   result_col109[55] <= result_col109[54];
   result_col109[56] <= result_col109[55];
   result_col109[57] <= result_col109[56];

   result_col110[1] <= data_out_4_110;
   result_col110[2] <= result_col110[1];
   result_col110[3] <= result_col110[2];
   result_col110[4] <= result_col110[3];
   result_col110[5] <= result_col110[4];
   result_col110[6] <= result_col110[5];
   result_col110[7] <= result_col110[6];
   result_col110[8] <= result_col110[7];
   result_col110[9] <= result_col110[8];
   result_col110[10] <= result_col110[9];
   result_col110[11] <= result_col110[10];
   result_col110[12] <= result_col110[11];
   result_col110[13] <= result_col110[12];
   result_col110[14] <= result_col110[13];
   result_col110[15] <= result_col110[14];
   result_col110[16] <= result_col110[15];
   result_col110[17] <= result_col110[16];
   result_col110[18] <= result_col110[17];
   result_col110[19] <= result_col110[18];
   result_col110[20] <= result_col110[19];
   result_col110[21] <= result_col110[20];
   result_col110[22] <= result_col110[21];
   result_col110[23] <= result_col110[22];
   result_col110[24] <= result_col110[23];
   result_col110[25] <= result_col110[24];
   result_col110[26] <= result_col110[25];
   result_col110[27] <= result_col110[26];
   result_col110[28] <= result_col110[27];
   result_col110[29] <= result_col110[28];
   result_col110[30] <= result_col110[29];
   result_col110[31] <= result_col110[30];
   result_col110[32] <= result_col110[31];
   result_col110[33] <= result_col110[32];
   result_col110[34] <= result_col110[33];
   result_col110[35] <= result_col110[34];
   result_col110[36] <= result_col110[35];
   result_col110[37] <= result_col110[36];
   result_col110[38] <= result_col110[37];
   result_col110[39] <= result_col110[38];
   result_col110[40] <= result_col110[39];
   result_col110[41] <= result_col110[40];
   result_col110[42] <= result_col110[41];
   result_col110[43] <= result_col110[42];
   result_col110[44] <= result_col110[43];
   result_col110[45] <= result_col110[44];
   result_col110[46] <= result_col110[45];
   result_col110[47] <= result_col110[46];
   result_col110[48] <= result_col110[47];
   result_col110[49] <= result_col110[48];
   result_col110[50] <= result_col110[49];
   result_col110[51] <= result_col110[50];
   result_col110[52] <= result_col110[51];
   result_col110[53] <= result_col110[52];
   result_col110[54] <= result_col110[53];
   result_col110[55] <= result_col110[54];
   result_col110[56] <= result_col110[55];

   result_col111[1] <= data_out_4_111;
   result_col111[2] <= result_col111[1];
   result_col111[3] <= result_col111[2];
   result_col111[4] <= result_col111[3];
   result_col111[5] <= result_col111[4];
   result_col111[6] <= result_col111[5];
   result_col111[7] <= result_col111[6];
   result_col111[8] <= result_col111[7];
   result_col111[9] <= result_col111[8];
   result_col111[10] <= result_col111[9];
   result_col111[11] <= result_col111[10];
   result_col111[12] <= result_col111[11];
   result_col111[13] <= result_col111[12];
   result_col111[14] <= result_col111[13];
   result_col111[15] <= result_col111[14];
   result_col111[16] <= result_col111[15];
   result_col111[17] <= result_col111[16];
   result_col111[18] <= result_col111[17];
   result_col111[19] <= result_col111[18];
   result_col111[20] <= result_col111[19];
   result_col111[21] <= result_col111[20];
   result_col111[22] <= result_col111[21];
   result_col111[23] <= result_col111[22];
   result_col111[24] <= result_col111[23];
   result_col111[25] <= result_col111[24];
   result_col111[26] <= result_col111[25];
   result_col111[27] <= result_col111[26];
   result_col111[28] <= result_col111[27];
   result_col111[29] <= result_col111[28];
   result_col111[30] <= result_col111[29];
   result_col111[31] <= result_col111[30];
   result_col111[32] <= result_col111[31];
   result_col111[33] <= result_col111[32];
   result_col111[34] <= result_col111[33];
   result_col111[35] <= result_col111[34];
   result_col111[36] <= result_col111[35];
   result_col111[37] <= result_col111[36];
   result_col111[38] <= result_col111[37];
   result_col111[39] <= result_col111[38];
   result_col111[40] <= result_col111[39];
   result_col111[41] <= result_col111[40];
   result_col111[42] <= result_col111[41];
   result_col111[43] <= result_col111[42];
   result_col111[44] <= result_col111[43];
   result_col111[45] <= result_col111[44];
   result_col111[46] <= result_col111[45];
   result_col111[47] <= result_col111[46];
   result_col111[48] <= result_col111[47];
   result_col111[49] <= result_col111[48];
   result_col111[50] <= result_col111[49];
   result_col111[51] <= result_col111[50];
   result_col111[52] <= result_col111[51];
   result_col111[53] <= result_col111[52];
   result_col111[54] <= result_col111[53];
   result_col111[55] <= result_col111[54];

   result_col112[1] <= data_out_4_112;
   result_col112[2] <= result_col112[1];
   result_col112[3] <= result_col112[2];
   result_col112[4] <= result_col112[3];
   result_col112[5] <= result_col112[4];
   result_col112[6] <= result_col112[5];
   result_col112[7] <= result_col112[6];
   result_col112[8] <= result_col112[7];
   result_col112[9] <= result_col112[8];
   result_col112[10] <= result_col112[9];
   result_col112[11] <= result_col112[10];
   result_col112[12] <= result_col112[11];
   result_col112[13] <= result_col112[12];
   result_col112[14] <= result_col112[13];
   result_col112[15] <= result_col112[14];
   result_col112[16] <= result_col112[15];
   result_col112[17] <= result_col112[16];
   result_col112[18] <= result_col112[17];
   result_col112[19] <= result_col112[18];
   result_col112[20] <= result_col112[19];
   result_col112[21] <= result_col112[20];
   result_col112[22] <= result_col112[21];
   result_col112[23] <= result_col112[22];
   result_col112[24] <= result_col112[23];
   result_col112[25] <= result_col112[24];
   result_col112[26] <= result_col112[25];
   result_col112[27] <= result_col112[26];
   result_col112[28] <= result_col112[27];
   result_col112[29] <= result_col112[28];
   result_col112[30] <= result_col112[29];
   result_col112[31] <= result_col112[30];
   result_col112[32] <= result_col112[31];
   result_col112[33] <= result_col112[32];
   result_col112[34] <= result_col112[33];
   result_col112[35] <= result_col112[34];
   result_col112[36] <= result_col112[35];
   result_col112[37] <= result_col112[36];
   result_col112[38] <= result_col112[37];
   result_col112[39] <= result_col112[38];
   result_col112[40] <= result_col112[39];
   result_col112[41] <= result_col112[40];
   result_col112[42] <= result_col112[41];
   result_col112[43] <= result_col112[42];
   result_col112[44] <= result_col112[43];
   result_col112[45] <= result_col112[44];
   result_col112[46] <= result_col112[45];
   result_col112[47] <= result_col112[46];
   result_col112[48] <= result_col112[47];
   result_col112[49] <= result_col112[48];
   result_col112[50] <= result_col112[49];
   result_col112[51] <= result_col112[50];
   result_col112[52] <= result_col112[51];
   result_col112[53] <= result_col112[52];
   result_col112[54] <= result_col112[53];

   result_col113[1] <= data_out_4_113;
   result_col113[2] <= result_col113[1];
   result_col113[3] <= result_col113[2];
   result_col113[4] <= result_col113[3];
   result_col113[5] <= result_col113[4];
   result_col113[6] <= result_col113[5];
   result_col113[7] <= result_col113[6];
   result_col113[8] <= result_col113[7];
   result_col113[9] <= result_col113[8];
   result_col113[10] <= result_col113[9];
   result_col113[11] <= result_col113[10];
   result_col113[12] <= result_col113[11];
   result_col113[13] <= result_col113[12];
   result_col113[14] <= result_col113[13];
   result_col113[15] <= result_col113[14];
   result_col113[16] <= result_col113[15];
   result_col113[17] <= result_col113[16];
   result_col113[18] <= result_col113[17];
   result_col113[19] <= result_col113[18];
   result_col113[20] <= result_col113[19];
   result_col113[21] <= result_col113[20];
   result_col113[22] <= result_col113[21];
   result_col113[23] <= result_col113[22];
   result_col113[24] <= result_col113[23];
   result_col113[25] <= result_col113[24];
   result_col113[26] <= result_col113[25];
   result_col113[27] <= result_col113[26];
   result_col113[28] <= result_col113[27];
   result_col113[29] <= result_col113[28];
   result_col113[30] <= result_col113[29];
   result_col113[31] <= result_col113[30];
   result_col113[32] <= result_col113[31];
   result_col113[33] <= result_col113[32];
   result_col113[34] <= result_col113[33];
   result_col113[35] <= result_col113[34];
   result_col113[36] <= result_col113[35];
   result_col113[37] <= result_col113[36];
   result_col113[38] <= result_col113[37];
   result_col113[39] <= result_col113[38];
   result_col113[40] <= result_col113[39];
   result_col113[41] <= result_col113[40];
   result_col113[42] <= result_col113[41];
   result_col113[43] <= result_col113[42];
   result_col113[44] <= result_col113[43];
   result_col113[45] <= result_col113[44];
   result_col113[46] <= result_col113[45];
   result_col113[47] <= result_col113[46];
   result_col113[48] <= result_col113[47];
   result_col113[49] <= result_col113[48];
   result_col113[50] <= result_col113[49];
   result_col113[51] <= result_col113[50];
   result_col113[52] <= result_col113[51];
   result_col113[53] <= result_col113[52];

   result_col114[1] <= data_out_4_114;
   result_col114[2] <= result_col114[1];
   result_col114[3] <= result_col114[2];
   result_col114[4] <= result_col114[3];
   result_col114[5] <= result_col114[4];
   result_col114[6] <= result_col114[5];
   result_col114[7] <= result_col114[6];
   result_col114[8] <= result_col114[7];
   result_col114[9] <= result_col114[8];
   result_col114[10] <= result_col114[9];
   result_col114[11] <= result_col114[10];
   result_col114[12] <= result_col114[11];
   result_col114[13] <= result_col114[12];
   result_col114[14] <= result_col114[13];
   result_col114[15] <= result_col114[14];
   result_col114[16] <= result_col114[15];
   result_col114[17] <= result_col114[16];
   result_col114[18] <= result_col114[17];
   result_col114[19] <= result_col114[18];
   result_col114[20] <= result_col114[19];
   result_col114[21] <= result_col114[20];
   result_col114[22] <= result_col114[21];
   result_col114[23] <= result_col114[22];
   result_col114[24] <= result_col114[23];
   result_col114[25] <= result_col114[24];
   result_col114[26] <= result_col114[25];
   result_col114[27] <= result_col114[26];
   result_col114[28] <= result_col114[27];
   result_col114[29] <= result_col114[28];
   result_col114[30] <= result_col114[29];
   result_col114[31] <= result_col114[30];
   result_col114[32] <= result_col114[31];
   result_col114[33] <= result_col114[32];
   result_col114[34] <= result_col114[33];
   result_col114[35] <= result_col114[34];
   result_col114[36] <= result_col114[35];
   result_col114[37] <= result_col114[36];
   result_col114[38] <= result_col114[37];
   result_col114[39] <= result_col114[38];
   result_col114[40] <= result_col114[39];
   result_col114[41] <= result_col114[40];
   result_col114[42] <= result_col114[41];
   result_col114[43] <= result_col114[42];
   result_col114[44] <= result_col114[43];
   result_col114[45] <= result_col114[44];
   result_col114[46] <= result_col114[45];
   result_col114[47] <= result_col114[46];
   result_col114[48] <= result_col114[47];
   result_col114[49] <= result_col114[48];
   result_col114[50] <= result_col114[49];
   result_col114[51] <= result_col114[50];
   result_col114[52] <= result_col114[51];

   result_col115[1] <= data_out_4_115;
   result_col115[2] <= result_col115[1];
   result_col115[3] <= result_col115[2];
   result_col115[4] <= result_col115[3];
   result_col115[5] <= result_col115[4];
   result_col115[6] <= result_col115[5];
   result_col115[7] <= result_col115[6];
   result_col115[8] <= result_col115[7];
   result_col115[9] <= result_col115[8];
   result_col115[10] <= result_col115[9];
   result_col115[11] <= result_col115[10];
   result_col115[12] <= result_col115[11];
   result_col115[13] <= result_col115[12];
   result_col115[14] <= result_col115[13];
   result_col115[15] <= result_col115[14];
   result_col115[16] <= result_col115[15];
   result_col115[17] <= result_col115[16];
   result_col115[18] <= result_col115[17];
   result_col115[19] <= result_col115[18];
   result_col115[20] <= result_col115[19];
   result_col115[21] <= result_col115[20];
   result_col115[22] <= result_col115[21];
   result_col115[23] <= result_col115[22];
   result_col115[24] <= result_col115[23];
   result_col115[25] <= result_col115[24];
   result_col115[26] <= result_col115[25];
   result_col115[27] <= result_col115[26];
   result_col115[28] <= result_col115[27];
   result_col115[29] <= result_col115[28];
   result_col115[30] <= result_col115[29];
   result_col115[31] <= result_col115[30];
   result_col115[32] <= result_col115[31];
   result_col115[33] <= result_col115[32];
   result_col115[34] <= result_col115[33];
   result_col115[35] <= result_col115[34];
   result_col115[36] <= result_col115[35];
   result_col115[37] <= result_col115[36];
   result_col115[38] <= result_col115[37];
   result_col115[39] <= result_col115[38];
   result_col115[40] <= result_col115[39];
   result_col115[41] <= result_col115[40];
   result_col115[42] <= result_col115[41];
   result_col115[43] <= result_col115[42];
   result_col115[44] <= result_col115[43];
   result_col115[45] <= result_col115[44];
   result_col115[46] <= result_col115[45];
   result_col115[47] <= result_col115[46];
   result_col115[48] <= result_col115[47];
   result_col115[49] <= result_col115[48];
   result_col115[50] <= result_col115[49];
   result_col115[51] <= result_col115[50];

   result_col116[1] <= data_out_4_116;
   result_col116[2] <= result_col116[1];
   result_col116[3] <= result_col116[2];
   result_col116[4] <= result_col116[3];
   result_col116[5] <= result_col116[4];
   result_col116[6] <= result_col116[5];
   result_col116[7] <= result_col116[6];
   result_col116[8] <= result_col116[7];
   result_col116[9] <= result_col116[8];
   result_col116[10] <= result_col116[9];
   result_col116[11] <= result_col116[10];
   result_col116[12] <= result_col116[11];
   result_col116[13] <= result_col116[12];
   result_col116[14] <= result_col116[13];
   result_col116[15] <= result_col116[14];
   result_col116[16] <= result_col116[15];
   result_col116[17] <= result_col116[16];
   result_col116[18] <= result_col116[17];
   result_col116[19] <= result_col116[18];
   result_col116[20] <= result_col116[19];
   result_col116[21] <= result_col116[20];
   result_col116[22] <= result_col116[21];
   result_col116[23] <= result_col116[22];
   result_col116[24] <= result_col116[23];
   result_col116[25] <= result_col116[24];
   result_col116[26] <= result_col116[25];
   result_col116[27] <= result_col116[26];
   result_col116[28] <= result_col116[27];
   result_col116[29] <= result_col116[28];
   result_col116[30] <= result_col116[29];
   result_col116[31] <= result_col116[30];
   result_col116[32] <= result_col116[31];
   result_col116[33] <= result_col116[32];
   result_col116[34] <= result_col116[33];
   result_col116[35] <= result_col116[34];
   result_col116[36] <= result_col116[35];
   result_col116[37] <= result_col116[36];
   result_col116[38] <= result_col116[37];
   result_col116[39] <= result_col116[38];
   result_col116[40] <= result_col116[39];
   result_col116[41] <= result_col116[40];
   result_col116[42] <= result_col116[41];
   result_col116[43] <= result_col116[42];
   result_col116[44] <= result_col116[43];
   result_col116[45] <= result_col116[44];
   result_col116[46] <= result_col116[45];
   result_col116[47] <= result_col116[46];
   result_col116[48] <= result_col116[47];
   result_col116[49] <= result_col116[48];
   result_col116[50] <= result_col116[49];

   result_col117[1] <= data_out_4_117;
   result_col117[2] <= result_col117[1];
   result_col117[3] <= result_col117[2];
   result_col117[4] <= result_col117[3];
   result_col117[5] <= result_col117[4];
   result_col117[6] <= result_col117[5];
   result_col117[7] <= result_col117[6];
   result_col117[8] <= result_col117[7];
   result_col117[9] <= result_col117[8];
   result_col117[10] <= result_col117[9];
   result_col117[11] <= result_col117[10];
   result_col117[12] <= result_col117[11];
   result_col117[13] <= result_col117[12];
   result_col117[14] <= result_col117[13];
   result_col117[15] <= result_col117[14];
   result_col117[16] <= result_col117[15];
   result_col117[17] <= result_col117[16];
   result_col117[18] <= result_col117[17];
   result_col117[19] <= result_col117[18];
   result_col117[20] <= result_col117[19];
   result_col117[21] <= result_col117[20];
   result_col117[22] <= result_col117[21];
   result_col117[23] <= result_col117[22];
   result_col117[24] <= result_col117[23];
   result_col117[25] <= result_col117[24];
   result_col117[26] <= result_col117[25];
   result_col117[27] <= result_col117[26];
   result_col117[28] <= result_col117[27];
   result_col117[29] <= result_col117[28];
   result_col117[30] <= result_col117[29];
   result_col117[31] <= result_col117[30];
   result_col117[32] <= result_col117[31];
   result_col117[33] <= result_col117[32];
   result_col117[34] <= result_col117[33];
   result_col117[35] <= result_col117[34];
   result_col117[36] <= result_col117[35];
   result_col117[37] <= result_col117[36];
   result_col117[38] <= result_col117[37];
   result_col117[39] <= result_col117[38];
   result_col117[40] <= result_col117[39];
   result_col117[41] <= result_col117[40];
   result_col117[42] <= result_col117[41];
   result_col117[43] <= result_col117[42];
   result_col117[44] <= result_col117[43];
   result_col117[45] <= result_col117[44];
   result_col117[46] <= result_col117[45];
   result_col117[47] <= result_col117[46];
   result_col117[48] <= result_col117[47];
   result_col117[49] <= result_col117[48];

   result_col118[1] <= data_out_4_118;
   result_col118[2] <= result_col118[1];
   result_col118[3] <= result_col118[2];
   result_col118[4] <= result_col118[3];
   result_col118[5] <= result_col118[4];
   result_col118[6] <= result_col118[5];
   result_col118[7] <= result_col118[6];
   result_col118[8] <= result_col118[7];
   result_col118[9] <= result_col118[8];
   result_col118[10] <= result_col118[9];
   result_col118[11] <= result_col118[10];
   result_col118[12] <= result_col118[11];
   result_col118[13] <= result_col118[12];
   result_col118[14] <= result_col118[13];
   result_col118[15] <= result_col118[14];
   result_col118[16] <= result_col118[15];
   result_col118[17] <= result_col118[16];
   result_col118[18] <= result_col118[17];
   result_col118[19] <= result_col118[18];
   result_col118[20] <= result_col118[19];
   result_col118[21] <= result_col118[20];
   result_col118[22] <= result_col118[21];
   result_col118[23] <= result_col118[22];
   result_col118[24] <= result_col118[23];
   result_col118[25] <= result_col118[24];
   result_col118[26] <= result_col118[25];
   result_col118[27] <= result_col118[26];
   result_col118[28] <= result_col118[27];
   result_col118[29] <= result_col118[28];
   result_col118[30] <= result_col118[29];
   result_col118[31] <= result_col118[30];
   result_col118[32] <= result_col118[31];
   result_col118[33] <= result_col118[32];
   result_col118[34] <= result_col118[33];
   result_col118[35] <= result_col118[34];
   result_col118[36] <= result_col118[35];
   result_col118[37] <= result_col118[36];
   result_col118[38] <= result_col118[37];
   result_col118[39] <= result_col118[38];
   result_col118[40] <= result_col118[39];
   result_col118[41] <= result_col118[40];
   result_col118[42] <= result_col118[41];
   result_col118[43] <= result_col118[42];
   result_col118[44] <= result_col118[43];
   result_col118[45] <= result_col118[44];
   result_col118[46] <= result_col118[45];
   result_col118[47] <= result_col118[46];
   result_col118[48] <= result_col118[47];

   result_col119[1] <= data_out_4_119;
   result_col119[2] <= result_col119[1];
   result_col119[3] <= result_col119[2];
   result_col119[4] <= result_col119[3];
   result_col119[5] <= result_col119[4];
   result_col119[6] <= result_col119[5];
   result_col119[7] <= result_col119[6];
   result_col119[8] <= result_col119[7];
   result_col119[9] <= result_col119[8];
   result_col119[10] <= result_col119[9];
   result_col119[11] <= result_col119[10];
   result_col119[12] <= result_col119[11];
   result_col119[13] <= result_col119[12];
   result_col119[14] <= result_col119[13];
   result_col119[15] <= result_col119[14];
   result_col119[16] <= result_col119[15];
   result_col119[17] <= result_col119[16];
   result_col119[18] <= result_col119[17];
   result_col119[19] <= result_col119[18];
   result_col119[20] <= result_col119[19];
   result_col119[21] <= result_col119[20];
   result_col119[22] <= result_col119[21];
   result_col119[23] <= result_col119[22];
   result_col119[24] <= result_col119[23];
   result_col119[25] <= result_col119[24];
   result_col119[26] <= result_col119[25];
   result_col119[27] <= result_col119[26];
   result_col119[28] <= result_col119[27];
   result_col119[29] <= result_col119[28];
   result_col119[30] <= result_col119[29];
   result_col119[31] <= result_col119[30];
   result_col119[32] <= result_col119[31];
   result_col119[33] <= result_col119[32];
   result_col119[34] <= result_col119[33];
   result_col119[35] <= result_col119[34];
   result_col119[36] <= result_col119[35];
   result_col119[37] <= result_col119[36];
   result_col119[38] <= result_col119[37];
   result_col119[39] <= result_col119[38];
   result_col119[40] <= result_col119[39];
   result_col119[41] <= result_col119[40];
   result_col119[42] <= result_col119[41];
   result_col119[43] <= result_col119[42];
   result_col119[44] <= result_col119[43];
   result_col119[45] <= result_col119[44];
   result_col119[46] <= result_col119[45];
   result_col119[47] <= result_col119[46];

   result_col120[1] <= data_out_4_120;
   result_col120[2] <= result_col120[1];
   result_col120[3] <= result_col120[2];
   result_col120[4] <= result_col120[3];
   result_col120[5] <= result_col120[4];
   result_col120[6] <= result_col120[5];
   result_col120[7] <= result_col120[6];
   result_col120[8] <= result_col120[7];
   result_col120[9] <= result_col120[8];
   result_col120[10] <= result_col120[9];
   result_col120[11] <= result_col120[10];
   result_col120[12] <= result_col120[11];
   result_col120[13] <= result_col120[12];
   result_col120[14] <= result_col120[13];
   result_col120[15] <= result_col120[14];
   result_col120[16] <= result_col120[15];
   result_col120[17] <= result_col120[16];
   result_col120[18] <= result_col120[17];
   result_col120[19] <= result_col120[18];
   result_col120[20] <= result_col120[19];
   result_col120[21] <= result_col120[20];
   result_col120[22] <= result_col120[21];
   result_col120[23] <= result_col120[22];
   result_col120[24] <= result_col120[23];
   result_col120[25] <= result_col120[24];
   result_col120[26] <= result_col120[25];
   result_col120[27] <= result_col120[26];
   result_col120[28] <= result_col120[27];
   result_col120[29] <= result_col120[28];
   result_col120[30] <= result_col120[29];
   result_col120[31] <= result_col120[30];
   result_col120[32] <= result_col120[31];
   result_col120[33] <= result_col120[32];
   result_col120[34] <= result_col120[33];
   result_col120[35] <= result_col120[34];
   result_col120[36] <= result_col120[35];
   result_col120[37] <= result_col120[36];
   result_col120[38] <= result_col120[37];
   result_col120[39] <= result_col120[38];
   result_col120[40] <= result_col120[39];
   result_col120[41] <= result_col120[40];
   result_col120[42] <= result_col120[41];
   result_col120[43] <= result_col120[42];
   result_col120[44] <= result_col120[43];
   result_col120[45] <= result_col120[44];
   result_col120[46] <= result_col120[45];

   result_col121[1] <= data_out_4_121;
   result_col121[2] <= result_col121[1];
   result_col121[3] <= result_col121[2];
   result_col121[4] <= result_col121[3];
   result_col121[5] <= result_col121[4];
   result_col121[6] <= result_col121[5];
   result_col121[7] <= result_col121[6];
   result_col121[8] <= result_col121[7];
   result_col121[9] <= result_col121[8];
   result_col121[10] <= result_col121[9];
   result_col121[11] <= result_col121[10];
   result_col121[12] <= result_col121[11];
   result_col121[13] <= result_col121[12];
   result_col121[14] <= result_col121[13];
   result_col121[15] <= result_col121[14];
   result_col121[16] <= result_col121[15];
   result_col121[17] <= result_col121[16];
   result_col121[18] <= result_col121[17];
   result_col121[19] <= result_col121[18];
   result_col121[20] <= result_col121[19];
   result_col121[21] <= result_col121[20];
   result_col121[22] <= result_col121[21];
   result_col121[23] <= result_col121[22];
   result_col121[24] <= result_col121[23];
   result_col121[25] <= result_col121[24];
   result_col121[26] <= result_col121[25];
   result_col121[27] <= result_col121[26];
   result_col121[28] <= result_col121[27];
   result_col121[29] <= result_col121[28];
   result_col121[30] <= result_col121[29];
   result_col121[31] <= result_col121[30];
   result_col121[32] <= result_col121[31];
   result_col121[33] <= result_col121[32];
   result_col121[34] <= result_col121[33];
   result_col121[35] <= result_col121[34];
   result_col121[36] <= result_col121[35];
   result_col121[37] <= result_col121[36];
   result_col121[38] <= result_col121[37];
   result_col121[39] <= result_col121[38];
   result_col121[40] <= result_col121[39];
   result_col121[41] <= result_col121[40];
   result_col121[42] <= result_col121[41];
   result_col121[43] <= result_col121[42];
   result_col121[44] <= result_col121[43];
   result_col121[45] <= result_col121[44];

   result_col122[1] <= data_out_4_122;
   result_col122[2] <= result_col122[1];
   result_col122[3] <= result_col122[2];
   result_col122[4] <= result_col122[3];
   result_col122[5] <= result_col122[4];
   result_col122[6] <= result_col122[5];
   result_col122[7] <= result_col122[6];
   result_col122[8] <= result_col122[7];
   result_col122[9] <= result_col122[8];
   result_col122[10] <= result_col122[9];
   result_col122[11] <= result_col122[10];
   result_col122[12] <= result_col122[11];
   result_col122[13] <= result_col122[12];
   result_col122[14] <= result_col122[13];
   result_col122[15] <= result_col122[14];
   result_col122[16] <= result_col122[15];
   result_col122[17] <= result_col122[16];
   result_col122[18] <= result_col122[17];
   result_col122[19] <= result_col122[18];
   result_col122[20] <= result_col122[19];
   result_col122[21] <= result_col122[20];
   result_col122[22] <= result_col122[21];
   result_col122[23] <= result_col122[22];
   result_col122[24] <= result_col122[23];
   result_col122[25] <= result_col122[24];
   result_col122[26] <= result_col122[25];
   result_col122[27] <= result_col122[26];
   result_col122[28] <= result_col122[27];
   result_col122[29] <= result_col122[28];
   result_col122[30] <= result_col122[29];
   result_col122[31] <= result_col122[30];
   result_col122[32] <= result_col122[31];
   result_col122[33] <= result_col122[32];
   result_col122[34] <= result_col122[33];
   result_col122[35] <= result_col122[34];
   result_col122[36] <= result_col122[35];
   result_col122[37] <= result_col122[36];
   result_col122[38] <= result_col122[37];
   result_col122[39] <= result_col122[38];
   result_col122[40] <= result_col122[39];
   result_col122[41] <= result_col122[40];
   result_col122[42] <= result_col122[41];
   result_col122[43] <= result_col122[42];
   result_col122[44] <= result_col122[43];

   result_col123[1] <= data_out_4_123;
   result_col123[2] <= result_col123[1];
   result_col123[3] <= result_col123[2];
   result_col123[4] <= result_col123[3];
   result_col123[5] <= result_col123[4];
   result_col123[6] <= result_col123[5];
   result_col123[7] <= result_col123[6];
   result_col123[8] <= result_col123[7];
   result_col123[9] <= result_col123[8];
   result_col123[10] <= result_col123[9];
   result_col123[11] <= result_col123[10];
   result_col123[12] <= result_col123[11];
   result_col123[13] <= result_col123[12];
   result_col123[14] <= result_col123[13];
   result_col123[15] <= result_col123[14];
   result_col123[16] <= result_col123[15];
   result_col123[17] <= result_col123[16];
   result_col123[18] <= result_col123[17];
   result_col123[19] <= result_col123[18];
   result_col123[20] <= result_col123[19];
   result_col123[21] <= result_col123[20];
   result_col123[22] <= result_col123[21];
   result_col123[23] <= result_col123[22];
   result_col123[24] <= result_col123[23];
   result_col123[25] <= result_col123[24];
   result_col123[26] <= result_col123[25];
   result_col123[27] <= result_col123[26];
   result_col123[28] <= result_col123[27];
   result_col123[29] <= result_col123[28];
   result_col123[30] <= result_col123[29];
   result_col123[31] <= result_col123[30];
   result_col123[32] <= result_col123[31];
   result_col123[33] <= result_col123[32];
   result_col123[34] <= result_col123[33];
   result_col123[35] <= result_col123[34];
   result_col123[36] <= result_col123[35];
   result_col123[37] <= result_col123[36];
   result_col123[38] <= result_col123[37];
   result_col123[39] <= result_col123[38];
   result_col123[40] <= result_col123[39];
   result_col123[41] <= result_col123[40];
   result_col123[42] <= result_col123[41];
   result_col123[43] <= result_col123[42];

   result_col124[1] <= data_out_4_124;
   result_col124[2] <= result_col124[1];
   result_col124[3] <= result_col124[2];
   result_col124[4] <= result_col124[3];
   result_col124[5] <= result_col124[4];
   result_col124[6] <= result_col124[5];
   result_col124[7] <= result_col124[6];
   result_col124[8] <= result_col124[7];
   result_col124[9] <= result_col124[8];
   result_col124[10] <= result_col124[9];
   result_col124[11] <= result_col124[10];
   result_col124[12] <= result_col124[11];
   result_col124[13] <= result_col124[12];
   result_col124[14] <= result_col124[13];
   result_col124[15] <= result_col124[14];
   result_col124[16] <= result_col124[15];
   result_col124[17] <= result_col124[16];
   result_col124[18] <= result_col124[17];
   result_col124[19] <= result_col124[18];
   result_col124[20] <= result_col124[19];
   result_col124[21] <= result_col124[20];
   result_col124[22] <= result_col124[21];
   result_col124[23] <= result_col124[22];
   result_col124[24] <= result_col124[23];
   result_col124[25] <= result_col124[24];
   result_col124[26] <= result_col124[25];
   result_col124[27] <= result_col124[26];
   result_col124[28] <= result_col124[27];
   result_col124[29] <= result_col124[28];
   result_col124[30] <= result_col124[29];
   result_col124[31] <= result_col124[30];
   result_col124[32] <= result_col124[31];
   result_col124[33] <= result_col124[32];
   result_col124[34] <= result_col124[33];
   result_col124[35] <= result_col124[34];
   result_col124[36] <= result_col124[35];
   result_col124[37] <= result_col124[36];
   result_col124[38] <= result_col124[37];
   result_col124[39] <= result_col124[38];
   result_col124[40] <= result_col124[39];
   result_col124[41] <= result_col124[40];
   result_col124[42] <= result_col124[41];

   result_col125[1] <= data_out_4_125;
   result_col125[2] <= result_col125[1];
   result_col125[3] <= result_col125[2];
   result_col125[4] <= result_col125[3];
   result_col125[5] <= result_col125[4];
   result_col125[6] <= result_col125[5];
   result_col125[7] <= result_col125[6];
   result_col125[8] <= result_col125[7];
   result_col125[9] <= result_col125[8];
   result_col125[10] <= result_col125[9];
   result_col125[11] <= result_col125[10];
   result_col125[12] <= result_col125[11];
   result_col125[13] <= result_col125[12];
   result_col125[14] <= result_col125[13];
   result_col125[15] <= result_col125[14];
   result_col125[16] <= result_col125[15];
   result_col125[17] <= result_col125[16];
   result_col125[18] <= result_col125[17];
   result_col125[19] <= result_col125[18];
   result_col125[20] <= result_col125[19];
   result_col125[21] <= result_col125[20];
   result_col125[22] <= result_col125[21];
   result_col125[23] <= result_col125[22];
   result_col125[24] <= result_col125[23];
   result_col125[25] <= result_col125[24];
   result_col125[26] <= result_col125[25];
   result_col125[27] <= result_col125[26];
   result_col125[28] <= result_col125[27];
   result_col125[29] <= result_col125[28];
   result_col125[30] <= result_col125[29];
   result_col125[31] <= result_col125[30];
   result_col125[32] <= result_col125[31];
   result_col125[33] <= result_col125[32];
   result_col125[34] <= result_col125[33];
   result_col125[35] <= result_col125[34];
   result_col125[36] <= result_col125[35];
   result_col125[37] <= result_col125[36];
   result_col125[38] <= result_col125[37];
   result_col125[39] <= result_col125[38];
   result_col125[40] <= result_col125[39];
   result_col125[41] <= result_col125[40];

   result_col126[1] <= data_out_4_126;
   result_col126[2] <= result_col126[1];
   result_col126[3] <= result_col126[2];
   result_col126[4] <= result_col126[3];
   result_col126[5] <= result_col126[4];
   result_col126[6] <= result_col126[5];
   result_col126[7] <= result_col126[6];
   result_col126[8] <= result_col126[7];
   result_col126[9] <= result_col126[8];
   result_col126[10] <= result_col126[9];
   result_col126[11] <= result_col126[10];
   result_col126[12] <= result_col126[11];
   result_col126[13] <= result_col126[12];
   result_col126[14] <= result_col126[13];
   result_col126[15] <= result_col126[14];
   result_col126[16] <= result_col126[15];
   result_col126[17] <= result_col126[16];
   result_col126[18] <= result_col126[17];
   result_col126[19] <= result_col126[18];
   result_col126[20] <= result_col126[19];
   result_col126[21] <= result_col126[20];
   result_col126[22] <= result_col126[21];
   result_col126[23] <= result_col126[22];
   result_col126[24] <= result_col126[23];
   result_col126[25] <= result_col126[24];
   result_col126[26] <= result_col126[25];
   result_col126[27] <= result_col126[26];
   result_col126[28] <= result_col126[27];
   result_col126[29] <= result_col126[28];
   result_col126[30] <= result_col126[29];
   result_col126[31] <= result_col126[30];
   result_col126[32] <= result_col126[31];
   result_col126[33] <= result_col126[32];
   result_col126[34] <= result_col126[33];
   result_col126[35] <= result_col126[34];
   result_col126[36] <= result_col126[35];
   result_col126[37] <= result_col126[36];
   result_col126[38] <= result_col126[37];
   result_col126[39] <= result_col126[38];
   result_col126[40] <= result_col126[39];

   result_col127[1] <= data_out_4_127;
   result_col127[2] <= result_col127[1];
   result_col127[3] <= result_col127[2];
   result_col127[4] <= result_col127[3];
   result_col127[5] <= result_col127[4];
   result_col127[6] <= result_col127[5];
   result_col127[7] <= result_col127[6];
   result_col127[8] <= result_col127[7];
   result_col127[9] <= result_col127[8];
   result_col127[10] <= result_col127[9];
   result_col127[11] <= result_col127[10];
   result_col127[12] <= result_col127[11];
   result_col127[13] <= result_col127[12];
   result_col127[14] <= result_col127[13];
   result_col127[15] <= result_col127[14];
   result_col127[16] <= result_col127[15];
   result_col127[17] <= result_col127[16];
   result_col127[18] <= result_col127[17];
   result_col127[19] <= result_col127[18];
   result_col127[20] <= result_col127[19];
   result_col127[21] <= result_col127[20];
   result_col127[22] <= result_col127[21];
   result_col127[23] <= result_col127[22];
   result_col127[24] <= result_col127[23];
   result_col127[25] <= result_col127[24];
   result_col127[26] <= result_col127[25];
   result_col127[27] <= result_col127[26];
   result_col127[28] <= result_col127[27];
   result_col127[29] <= result_col127[28];
   result_col127[30] <= result_col127[29];
   result_col127[31] <= result_col127[30];
   result_col127[32] <= result_col127[31];
   result_col127[33] <= result_col127[32];
   result_col127[34] <= result_col127[33];
   result_col127[35] <= result_col127[34];
   result_col127[36] <= result_col127[35];
   result_col127[37] <= result_col127[36];
   result_col127[38] <= result_col127[37];
   result_col127[39] <= result_col127[38];

   result_col128[1] <= data_out_4_128;
   result_col128[2] <= result_col128[1];
   result_col128[3] <= result_col128[2];
   result_col128[4] <= result_col128[3];
   result_col128[5] <= result_col128[4];
   result_col128[6] <= result_col128[5];
   result_col128[7] <= result_col128[6];
   result_col128[8] <= result_col128[7];
   result_col128[9] <= result_col128[8];
   result_col128[10] <= result_col128[9];
   result_col128[11] <= result_col128[10];
   result_col128[12] <= result_col128[11];
   result_col128[13] <= result_col128[12];
   result_col128[14] <= result_col128[13];
   result_col128[15] <= result_col128[14];
   result_col128[16] <= result_col128[15];
   result_col128[17] <= result_col128[16];
   result_col128[18] <= result_col128[17];
   result_col128[19] <= result_col128[18];
   result_col128[20] <= result_col128[19];
   result_col128[21] <= result_col128[20];
   result_col128[22] <= result_col128[21];
   result_col128[23] <= result_col128[22];
   result_col128[24] <= result_col128[23];
   result_col128[25] <= result_col128[24];
   result_col128[26] <= result_col128[25];
   result_col128[27] <= result_col128[26];
   result_col128[28] <= result_col128[27];
   result_col128[29] <= result_col128[28];
   result_col128[30] <= result_col128[29];
   result_col128[31] <= result_col128[30];
   result_col128[32] <= result_col128[31];
   result_col128[33] <= result_col128[32];
   result_col128[34] <= result_col128[33];
   result_col128[35] <= result_col128[34];
   result_col128[36] <= result_col128[35];
   result_col128[37] <= result_col128[36];
   result_col128[38] <= result_col128[37];

   result_col129[1] <= data_out_4_129;
   result_col129[2] <= result_col129[1];
   result_col129[3] <= result_col129[2];
   result_col129[4] <= result_col129[3];
   result_col129[5] <= result_col129[4];
   result_col129[6] <= result_col129[5];
   result_col129[7] <= result_col129[6];
   result_col129[8] <= result_col129[7];
   result_col129[9] <= result_col129[8];
   result_col129[10] <= result_col129[9];
   result_col129[11] <= result_col129[10];
   result_col129[12] <= result_col129[11];
   result_col129[13] <= result_col129[12];
   result_col129[14] <= result_col129[13];
   result_col129[15] <= result_col129[14];
   result_col129[16] <= result_col129[15];
   result_col129[17] <= result_col129[16];
   result_col129[18] <= result_col129[17];
   result_col129[19] <= result_col129[18];
   result_col129[20] <= result_col129[19];
   result_col129[21] <= result_col129[20];
   result_col129[22] <= result_col129[21];
   result_col129[23] <= result_col129[22];
   result_col129[24] <= result_col129[23];
   result_col129[25] <= result_col129[24];
   result_col129[26] <= result_col129[25];
   result_col129[27] <= result_col129[26];
   result_col129[28] <= result_col129[27];
   result_col129[29] <= result_col129[28];
   result_col129[30] <= result_col129[29];
   result_col129[31] <= result_col129[30];
   result_col129[32] <= result_col129[31];
   result_col129[33] <= result_col129[32];
   result_col129[34] <= result_col129[33];
   result_col129[35] <= result_col129[34];
   result_col129[36] <= result_col129[35];
   result_col129[37] <= result_col129[36];

   result_col130[1] <= data_out_4_130;
   result_col130[2] <= result_col130[1];
   result_col130[3] <= result_col130[2];
   result_col130[4] <= result_col130[3];
   result_col130[5] <= result_col130[4];
   result_col130[6] <= result_col130[5];
   result_col130[7] <= result_col130[6];
   result_col130[8] <= result_col130[7];
   result_col130[9] <= result_col130[8];
   result_col130[10] <= result_col130[9];
   result_col130[11] <= result_col130[10];
   result_col130[12] <= result_col130[11];
   result_col130[13] <= result_col130[12];
   result_col130[14] <= result_col130[13];
   result_col130[15] <= result_col130[14];
   result_col130[16] <= result_col130[15];
   result_col130[17] <= result_col130[16];
   result_col130[18] <= result_col130[17];
   result_col130[19] <= result_col130[18];
   result_col130[20] <= result_col130[19];
   result_col130[21] <= result_col130[20];
   result_col130[22] <= result_col130[21];
   result_col130[23] <= result_col130[22];
   result_col130[24] <= result_col130[23];
   result_col130[25] <= result_col130[24];
   result_col130[26] <= result_col130[25];
   result_col130[27] <= result_col130[26];
   result_col130[28] <= result_col130[27];
   result_col130[29] <= result_col130[28];
   result_col130[30] <= result_col130[29];
   result_col130[31] <= result_col130[30];
   result_col130[32] <= result_col130[31];
   result_col130[33] <= result_col130[32];
   result_col130[34] <= result_col130[33];
   result_col130[35] <= result_col130[34];
   result_col130[36] <= result_col130[35];

   result_col131[1] <= data_out_4_131;
   result_col131[2] <= result_col131[1];
   result_col131[3] <= result_col131[2];
   result_col131[4] <= result_col131[3];
   result_col131[5] <= result_col131[4];
   result_col131[6] <= result_col131[5];
   result_col131[7] <= result_col131[6];
   result_col131[8] <= result_col131[7];
   result_col131[9] <= result_col131[8];
   result_col131[10] <= result_col131[9];
   result_col131[11] <= result_col131[10];
   result_col131[12] <= result_col131[11];
   result_col131[13] <= result_col131[12];
   result_col131[14] <= result_col131[13];
   result_col131[15] <= result_col131[14];
   result_col131[16] <= result_col131[15];
   result_col131[17] <= result_col131[16];
   result_col131[18] <= result_col131[17];
   result_col131[19] <= result_col131[18];
   result_col131[20] <= result_col131[19];
   result_col131[21] <= result_col131[20];
   result_col131[22] <= result_col131[21];
   result_col131[23] <= result_col131[22];
   result_col131[24] <= result_col131[23];
   result_col131[25] <= result_col131[24];
   result_col131[26] <= result_col131[25];
   result_col131[27] <= result_col131[26];
   result_col131[28] <= result_col131[27];
   result_col131[29] <= result_col131[28];
   result_col131[30] <= result_col131[29];
   result_col131[31] <= result_col131[30];
   result_col131[32] <= result_col131[31];
   result_col131[33] <= result_col131[32];
   result_col131[34] <= result_col131[33];
   result_col131[35] <= result_col131[34];

   result_col132[1] <= data_out_4_132;
   result_col132[2] <= result_col132[1];
   result_col132[3] <= result_col132[2];
   result_col132[4] <= result_col132[3];
   result_col132[5] <= result_col132[4];
   result_col132[6] <= result_col132[5];
   result_col132[7] <= result_col132[6];
   result_col132[8] <= result_col132[7];
   result_col132[9] <= result_col132[8];
   result_col132[10] <= result_col132[9];
   result_col132[11] <= result_col132[10];
   result_col132[12] <= result_col132[11];
   result_col132[13] <= result_col132[12];
   result_col132[14] <= result_col132[13];
   result_col132[15] <= result_col132[14];
   result_col132[16] <= result_col132[15];
   result_col132[17] <= result_col132[16];
   result_col132[18] <= result_col132[17];
   result_col132[19] <= result_col132[18];
   result_col132[20] <= result_col132[19];
   result_col132[21] <= result_col132[20];
   result_col132[22] <= result_col132[21];
   result_col132[23] <= result_col132[22];
   result_col132[24] <= result_col132[23];
   result_col132[25] <= result_col132[24];
   result_col132[26] <= result_col132[25];
   result_col132[27] <= result_col132[26];
   result_col132[28] <= result_col132[27];
   result_col132[29] <= result_col132[28];
   result_col132[30] <= result_col132[29];
   result_col132[31] <= result_col132[30];
   result_col132[32] <= result_col132[31];
   result_col132[33] <= result_col132[32];
   result_col132[34] <= result_col132[33];

   result_col133[1] <= data_out_4_133;
   result_col133[2] <= result_col133[1];
   result_col133[3] <= result_col133[2];
   result_col133[4] <= result_col133[3];
   result_col133[5] <= result_col133[4];
   result_col133[6] <= result_col133[5];
   result_col133[7] <= result_col133[6];
   result_col133[8] <= result_col133[7];
   result_col133[9] <= result_col133[8];
   result_col133[10] <= result_col133[9];
   result_col133[11] <= result_col133[10];
   result_col133[12] <= result_col133[11];
   result_col133[13] <= result_col133[12];
   result_col133[14] <= result_col133[13];
   result_col133[15] <= result_col133[14];
   result_col133[16] <= result_col133[15];
   result_col133[17] <= result_col133[16];
   result_col133[18] <= result_col133[17];
   result_col133[19] <= result_col133[18];
   result_col133[20] <= result_col133[19];
   result_col133[21] <= result_col133[20];
   result_col133[22] <= result_col133[21];
   result_col133[23] <= result_col133[22];
   result_col133[24] <= result_col133[23];
   result_col133[25] <= result_col133[24];
   result_col133[26] <= result_col133[25];
   result_col133[27] <= result_col133[26];
   result_col133[28] <= result_col133[27];
   result_col133[29] <= result_col133[28];
   result_col133[30] <= result_col133[29];
   result_col133[31] <= result_col133[30];
   result_col133[32] <= result_col133[31];
   result_col133[33] <= result_col133[32];

   result_col134[1] <= data_out_4_134;
   result_col134[2] <= result_col134[1];
   result_col134[3] <= result_col134[2];
   result_col134[4] <= result_col134[3];
   result_col134[5] <= result_col134[4];
   result_col134[6] <= result_col134[5];
   result_col134[7] <= result_col134[6];
   result_col134[8] <= result_col134[7];
   result_col134[9] <= result_col134[8];
   result_col134[10] <= result_col134[9];
   result_col134[11] <= result_col134[10];
   result_col134[12] <= result_col134[11];
   result_col134[13] <= result_col134[12];
   result_col134[14] <= result_col134[13];
   result_col134[15] <= result_col134[14];
   result_col134[16] <= result_col134[15];
   result_col134[17] <= result_col134[16];
   result_col134[18] <= result_col134[17];
   result_col134[19] <= result_col134[18];
   result_col134[20] <= result_col134[19];
   result_col134[21] <= result_col134[20];
   result_col134[22] <= result_col134[21];
   result_col134[23] <= result_col134[22];
   result_col134[24] <= result_col134[23];
   result_col134[25] <= result_col134[24];
   result_col134[26] <= result_col134[25];
   result_col134[27] <= result_col134[26];
   result_col134[28] <= result_col134[27];
   result_col134[29] <= result_col134[28];
   result_col134[30] <= result_col134[29];
   result_col134[31] <= result_col134[30];
   result_col134[32] <= result_col134[31];

   result_col135[1] <= data_out_4_135;
   result_col135[2] <= result_col135[1];
   result_col135[3] <= result_col135[2];
   result_col135[4] <= result_col135[3];
   result_col135[5] <= result_col135[4];
   result_col135[6] <= result_col135[5];
   result_col135[7] <= result_col135[6];
   result_col135[8] <= result_col135[7];
   result_col135[9] <= result_col135[8];
   result_col135[10] <= result_col135[9];
   result_col135[11] <= result_col135[10];
   result_col135[12] <= result_col135[11];
   result_col135[13] <= result_col135[12];
   result_col135[14] <= result_col135[13];
   result_col135[15] <= result_col135[14];
   result_col135[16] <= result_col135[15];
   result_col135[17] <= result_col135[16];
   result_col135[18] <= result_col135[17];
   result_col135[19] <= result_col135[18];
   result_col135[20] <= result_col135[19];
   result_col135[21] <= result_col135[20];
   result_col135[22] <= result_col135[21];
   result_col135[23] <= result_col135[22];
   result_col135[24] <= result_col135[23];
   result_col135[25] <= result_col135[24];
   result_col135[26] <= result_col135[25];
   result_col135[27] <= result_col135[26];
   result_col135[28] <= result_col135[27];
   result_col135[29] <= result_col135[28];
   result_col135[30] <= result_col135[29];
   result_col135[31] <= result_col135[30];

   result_col136[1] <= data_out_4_136;
   result_col136[2] <= result_col136[1];
   result_col136[3] <= result_col136[2];
   result_col136[4] <= result_col136[3];
   result_col136[5] <= result_col136[4];
   result_col136[6] <= result_col136[5];
   result_col136[7] <= result_col136[6];
   result_col136[8] <= result_col136[7];
   result_col136[9] <= result_col136[8];
   result_col136[10] <= result_col136[9];
   result_col136[11] <= result_col136[10];
   result_col136[12] <= result_col136[11];
   result_col136[13] <= result_col136[12];
   result_col136[14] <= result_col136[13];
   result_col136[15] <= result_col136[14];
   result_col136[16] <= result_col136[15];
   result_col136[17] <= result_col136[16];
   result_col136[18] <= result_col136[17];
   result_col136[19] <= result_col136[18];
   result_col136[20] <= result_col136[19];
   result_col136[21] <= result_col136[20];
   result_col136[22] <= result_col136[21];
   result_col136[23] <= result_col136[22];
   result_col136[24] <= result_col136[23];
   result_col136[25] <= result_col136[24];
   result_col136[26] <= result_col136[25];
   result_col136[27] <= result_col136[26];
   result_col136[28] <= result_col136[27];
   result_col136[29] <= result_col136[28];
   result_col136[30] <= result_col136[29];

   result_col137[1] <= data_out_4_137;
   result_col137[2] <= result_col137[1];
   result_col137[3] <= result_col137[2];
   result_col137[4] <= result_col137[3];
   result_col137[5] <= result_col137[4];
   result_col137[6] <= result_col137[5];
   result_col137[7] <= result_col137[6];
   result_col137[8] <= result_col137[7];
   result_col137[9] <= result_col137[8];
   result_col137[10] <= result_col137[9];
   result_col137[11] <= result_col137[10];
   result_col137[12] <= result_col137[11];
   result_col137[13] <= result_col137[12];
   result_col137[14] <= result_col137[13];
   result_col137[15] <= result_col137[14];
   result_col137[16] <= result_col137[15];
   result_col137[17] <= result_col137[16];
   result_col137[18] <= result_col137[17];
   result_col137[19] <= result_col137[18];
   result_col137[20] <= result_col137[19];
   result_col137[21] <= result_col137[20];
   result_col137[22] <= result_col137[21];
   result_col137[23] <= result_col137[22];
   result_col137[24] <= result_col137[23];
   result_col137[25] <= result_col137[24];
   result_col137[26] <= result_col137[25];
   result_col137[27] <= result_col137[26];
   result_col137[28] <= result_col137[27];
   result_col137[29] <= result_col137[28];

   result_col138[1] <= data_out_4_138;
   result_col138[2] <= result_col138[1];
   result_col138[3] <= result_col138[2];
   result_col138[4] <= result_col138[3];
   result_col138[5] <= result_col138[4];
   result_col138[6] <= result_col138[5];
   result_col138[7] <= result_col138[6];
   result_col138[8] <= result_col138[7];
   result_col138[9] <= result_col138[8];
   result_col138[10] <= result_col138[9];
   result_col138[11] <= result_col138[10];
   result_col138[12] <= result_col138[11];
   result_col138[13] <= result_col138[12];
   result_col138[14] <= result_col138[13];
   result_col138[15] <= result_col138[14];
   result_col138[16] <= result_col138[15];
   result_col138[17] <= result_col138[16];
   result_col138[18] <= result_col138[17];
   result_col138[19] <= result_col138[18];
   result_col138[20] <= result_col138[19];
   result_col138[21] <= result_col138[20];
   result_col138[22] <= result_col138[21];
   result_col138[23] <= result_col138[22];
   result_col138[24] <= result_col138[23];
   result_col138[25] <= result_col138[24];
   result_col138[26] <= result_col138[25];
   result_col138[27] <= result_col138[26];
   result_col138[28] <= result_col138[27];

   result_col139[1] <= data_out_4_139;
   result_col139[2] <= result_col139[1];
   result_col139[3] <= result_col139[2];
   result_col139[4] <= result_col139[3];
   result_col139[5] <= result_col139[4];
   result_col139[6] <= result_col139[5];
   result_col139[7] <= result_col139[6];
   result_col139[8] <= result_col139[7];
   result_col139[9] <= result_col139[8];
   result_col139[10] <= result_col139[9];
   result_col139[11] <= result_col139[10];
   result_col139[12] <= result_col139[11];
   result_col139[13] <= result_col139[12];
   result_col139[14] <= result_col139[13];
   result_col139[15] <= result_col139[14];
   result_col139[16] <= result_col139[15];
   result_col139[17] <= result_col139[16];
   result_col139[18] <= result_col139[17];
   result_col139[19] <= result_col139[18];
   result_col139[20] <= result_col139[19];
   result_col139[21] <= result_col139[20];
   result_col139[22] <= result_col139[21];
   result_col139[23] <= result_col139[22];
   result_col139[24] <= result_col139[23];
   result_col139[25] <= result_col139[24];
   result_col139[26] <= result_col139[25];
   result_col139[27] <= result_col139[26];

   result_col140[1] <= data_out_4_140;
   result_col140[2] <= result_col140[1];
   result_col140[3] <= result_col140[2];
   result_col140[4] <= result_col140[3];
   result_col140[5] <= result_col140[4];
   result_col140[6] <= result_col140[5];
   result_col140[7] <= result_col140[6];
   result_col140[8] <= result_col140[7];
   result_col140[9] <= result_col140[8];
   result_col140[10] <= result_col140[9];
   result_col140[11] <= result_col140[10];
   result_col140[12] <= result_col140[11];
   result_col140[13] <= result_col140[12];
   result_col140[14] <= result_col140[13];
   result_col140[15] <= result_col140[14];
   result_col140[16] <= result_col140[15];
   result_col140[17] <= result_col140[16];
   result_col140[18] <= result_col140[17];
   result_col140[19] <= result_col140[18];
   result_col140[20] <= result_col140[19];
   result_col140[21] <= result_col140[20];
   result_col140[22] <= result_col140[21];
   result_col140[23] <= result_col140[22];
   result_col140[24] <= result_col140[23];
   result_col140[25] <= result_col140[24];
   result_col140[26] <= result_col140[25];

   result_col141[1] <= data_out_4_141;
   result_col141[2] <= result_col141[1];
   result_col141[3] <= result_col141[2];
   result_col141[4] <= result_col141[3];
   result_col141[5] <= result_col141[4];
   result_col141[6] <= result_col141[5];
   result_col141[7] <= result_col141[6];
   result_col141[8] <= result_col141[7];
   result_col141[9] <= result_col141[8];
   result_col141[10] <= result_col141[9];
   result_col141[11] <= result_col141[10];
   result_col141[12] <= result_col141[11];
   result_col141[13] <= result_col141[12];
   result_col141[14] <= result_col141[13];
   result_col141[15] <= result_col141[14];
   result_col141[16] <= result_col141[15];
   result_col141[17] <= result_col141[16];
   result_col141[18] <= result_col141[17];
   result_col141[19] <= result_col141[18];
   result_col141[20] <= result_col141[19];
   result_col141[21] <= result_col141[20];
   result_col141[22] <= result_col141[21];
   result_col141[23] <= result_col141[22];
   result_col141[24] <= result_col141[23];
   result_col141[25] <= result_col141[24];

   result_col142[1] <= data_out_4_142;
   result_col142[2] <= result_col142[1];
   result_col142[3] <= result_col142[2];
   result_col142[4] <= result_col142[3];
   result_col142[5] <= result_col142[4];
   result_col142[6] <= result_col142[5];
   result_col142[7] <= result_col142[6];
   result_col142[8] <= result_col142[7];
   result_col142[9] <= result_col142[8];
   result_col142[10] <= result_col142[9];
   result_col142[11] <= result_col142[10];
   result_col142[12] <= result_col142[11];
   result_col142[13] <= result_col142[12];
   result_col142[14] <= result_col142[13];
   result_col142[15] <= result_col142[14];
   result_col142[16] <= result_col142[15];
   result_col142[17] <= result_col142[16];
   result_col142[18] <= result_col142[17];
   result_col142[19] <= result_col142[18];
   result_col142[20] <= result_col142[19];
   result_col142[21] <= result_col142[20];
   result_col142[22] <= result_col142[21];
   result_col142[23] <= result_col142[22];
   result_col142[24] <= result_col142[23];

   result_col143[1] <= data_out_4_143;
   result_col143[2] <= result_col143[1];
   result_col143[3] <= result_col143[2];
   result_col143[4] <= result_col143[3];
   result_col143[5] <= result_col143[4];
   result_col143[6] <= result_col143[5];
   result_col143[7] <= result_col143[6];
   result_col143[8] <= result_col143[7];
   result_col143[9] <= result_col143[8];
   result_col143[10] <= result_col143[9];
   result_col143[11] <= result_col143[10];
   result_col143[12] <= result_col143[11];
   result_col143[13] <= result_col143[12];
   result_col143[14] <= result_col143[13];
   result_col143[15] <= result_col143[14];
   result_col143[16] <= result_col143[15];
   result_col143[17] <= result_col143[16];
   result_col143[18] <= result_col143[17];
   result_col143[19] <= result_col143[18];
   result_col143[20] <= result_col143[19];
   result_col143[21] <= result_col143[20];
   result_col143[22] <= result_col143[21];
   result_col143[23] <= result_col143[22];

   result_col144[1] <= data_out_4_144;
   result_col144[2] <= result_col144[1];
   result_col144[3] <= result_col144[2];
   result_col144[4] <= result_col144[3];
   result_col144[5] <= result_col144[4];
   result_col144[6] <= result_col144[5];
   result_col144[7] <= result_col144[6];
   result_col144[8] <= result_col144[7];
   result_col144[9] <= result_col144[8];
   result_col144[10] <= result_col144[9];
   result_col144[11] <= result_col144[10];
   result_col144[12] <= result_col144[11];
   result_col144[13] <= result_col144[12];
   result_col144[14] <= result_col144[13];
   result_col144[15] <= result_col144[14];
   result_col144[16] <= result_col144[15];
   result_col144[17] <= result_col144[16];
   result_col144[18] <= result_col144[17];
   result_col144[19] <= result_col144[18];
   result_col144[20] <= result_col144[19];
   result_col144[21] <= result_col144[20];
   result_col144[22] <= result_col144[21];

   result_col145[1] <= data_out_4_145;
   result_col145[2] <= result_col145[1];
   result_col145[3] <= result_col145[2];
   result_col145[4] <= result_col145[3];
   result_col145[5] <= result_col145[4];
   result_col145[6] <= result_col145[5];
   result_col145[7] <= result_col145[6];
   result_col145[8] <= result_col145[7];
   result_col145[9] <= result_col145[8];
   result_col145[10] <= result_col145[9];
   result_col145[11] <= result_col145[10];
   result_col145[12] <= result_col145[11];
   result_col145[13] <= result_col145[12];
   result_col145[14] <= result_col145[13];
   result_col145[15] <= result_col145[14];
   result_col145[16] <= result_col145[15];
   result_col145[17] <= result_col145[16];
   result_col145[18] <= result_col145[17];
   result_col145[19] <= result_col145[18];
   result_col145[20] <= result_col145[19];
   result_col145[21] <= result_col145[20];

   result_col146[1] <= data_out_4_146;
   result_col146[2] <= result_col146[1];
   result_col146[3] <= result_col146[2];
   result_col146[4] <= result_col146[3];
   result_col146[5] <= result_col146[4];
   result_col146[6] <= result_col146[5];
   result_col146[7] <= result_col146[6];
   result_col146[8] <= result_col146[7];
   result_col146[9] <= result_col146[8];
   result_col146[10] <= result_col146[9];
   result_col146[11] <= result_col146[10];
   result_col146[12] <= result_col146[11];
   result_col146[13] <= result_col146[12];
   result_col146[14] <= result_col146[13];
   result_col146[15] <= result_col146[14];
   result_col146[16] <= result_col146[15];
   result_col146[17] <= result_col146[16];
   result_col146[18] <= result_col146[17];
   result_col146[19] <= result_col146[18];
   result_col146[20] <= result_col146[19];

   result_col147[1] <= data_out_4_147;
   result_col147[2] <= result_col147[1];
   result_col147[3] <= result_col147[2];
   result_col147[4] <= result_col147[3];
   result_col147[5] <= result_col147[4];
   result_col147[6] <= result_col147[5];
   result_col147[7] <= result_col147[6];
   result_col147[8] <= result_col147[7];
   result_col147[9] <= result_col147[8];
   result_col147[10] <= result_col147[9];
   result_col147[11] <= result_col147[10];
   result_col147[12] <= result_col147[11];
   result_col147[13] <= result_col147[12];
   result_col147[14] <= result_col147[13];
   result_col147[15] <= result_col147[14];
   result_col147[16] <= result_col147[15];
   result_col147[17] <= result_col147[16];
   result_col147[18] <= result_col147[17];
   result_col147[19] <= result_col147[18];

   result_col148[1] <= data_out_4_148;
   result_col148[2] <= result_col148[1];
   result_col148[3] <= result_col148[2];
   result_col148[4] <= result_col148[3];
   result_col148[5] <= result_col148[4];
   result_col148[6] <= result_col148[5];
   result_col148[7] <= result_col148[6];
   result_col148[8] <= result_col148[7];
   result_col148[9] <= result_col148[8];
   result_col148[10] <= result_col148[9];
   result_col148[11] <= result_col148[10];
   result_col148[12] <= result_col148[11];
   result_col148[13] <= result_col148[12];
   result_col148[14] <= result_col148[13];
   result_col148[15] <= result_col148[14];
   result_col148[16] <= result_col148[15];
   result_col148[17] <= result_col148[16];
   result_col148[18] <= result_col148[17];

   result_col149[1] <= data_out_4_149;
   result_col149[2] <= result_col149[1];
   result_col149[3] <= result_col149[2];
   result_col149[4] <= result_col149[3];
   result_col149[5] <= result_col149[4];
   result_col149[6] <= result_col149[5];
   result_col149[7] <= result_col149[6];
   result_col149[8] <= result_col149[7];
   result_col149[9] <= result_col149[8];
   result_col149[10] <= result_col149[9];
   result_col149[11] <= result_col149[10];
   result_col149[12] <= result_col149[11];
   result_col149[13] <= result_col149[12];
   result_col149[14] <= result_col149[13];
   result_col149[15] <= result_col149[14];
   result_col149[16] <= result_col149[15];
   result_col149[17] <= result_col149[16];

   result_col150[1] <= data_out_4_150;
   result_col150[2] <= result_col150[1];
   result_col150[3] <= result_col150[2];
   result_col150[4] <= result_col150[3];
   result_col150[5] <= result_col150[4];
   result_col150[6] <= result_col150[5];
   result_col150[7] <= result_col150[6];
   result_col150[8] <= result_col150[7];
   result_col150[9] <= result_col150[8];
   result_col150[10] <= result_col150[9];
   result_col150[11] <= result_col150[10];
   result_col150[12] <= result_col150[11];
   result_col150[13] <= result_col150[12];
   result_col150[14] <= result_col150[13];
   result_col150[15] <= result_col150[14];
   result_col150[16] <= result_col150[15];

   result_col151[1] <= data_out_4_151;
   result_col151[2] <= result_col151[1];
   result_col151[3] <= result_col151[2];
   result_col151[4] <= result_col151[3];
   result_col151[5] <= result_col151[4];
   result_col151[6] <= result_col151[5];
   result_col151[7] <= result_col151[6];
   result_col151[8] <= result_col151[7];
   result_col151[9] <= result_col151[8];
   result_col151[10] <= result_col151[9];
   result_col151[11] <= result_col151[10];
   result_col151[12] <= result_col151[11];
   result_col151[13] <= result_col151[12];
   result_col151[14] <= result_col151[13];
   result_col151[15] <= result_col151[14];

   result_col152[1] <= data_out_4_152;
   result_col152[2] <= result_col152[1];
   result_col152[3] <= result_col152[2];
   result_col152[4] <= result_col152[3];
   result_col152[5] <= result_col152[4];
   result_col152[6] <= result_col152[5];
   result_col152[7] <= result_col152[6];
   result_col152[8] <= result_col152[7];
   result_col152[9] <= result_col152[8];
   result_col152[10] <= result_col152[9];
   result_col152[11] <= result_col152[10];
   result_col152[12] <= result_col152[11];
   result_col152[13] <= result_col152[12];
   result_col152[14] <= result_col152[13];

   result_col153[1] <= data_out_4_153;
   result_col153[2] <= result_col153[1];
   result_col153[3] <= result_col153[2];
   result_col153[4] <= result_col153[3];
   result_col153[5] <= result_col153[4];
   result_col153[6] <= result_col153[5];
   result_col153[7] <= result_col153[6];
   result_col153[8] <= result_col153[7];
   result_col153[9] <= result_col153[8];
   result_col153[10] <= result_col153[9];
   result_col153[11] <= result_col153[10];
   result_col153[12] <= result_col153[11];
   result_col153[13] <= result_col153[12];

   result_col154[1] <= data_out_4_154;
   result_col154[2] <= result_col154[1];
   result_col154[3] <= result_col154[2];
   result_col154[4] <= result_col154[3];
   result_col154[5] <= result_col154[4];
   result_col154[6] <= result_col154[5];
   result_col154[7] <= result_col154[6];
   result_col154[8] <= result_col154[7];
   result_col154[9] <= result_col154[8];
   result_col154[10] <= result_col154[9];
   result_col154[11] <= result_col154[10];
   result_col154[12] <= result_col154[11];

   result_col155[1] <= data_out_4_155;
   result_col155[2] <= result_col155[1];
   result_col155[3] <= result_col155[2];
   result_col155[4] <= result_col155[3];
   result_col155[5] <= result_col155[4];
   result_col155[6] <= result_col155[5];
   result_col155[7] <= result_col155[6];
   result_col155[8] <= result_col155[7];
   result_col155[9] <= result_col155[8];
   result_col155[10] <= result_col155[9];
   result_col155[11] <= result_col155[10];

   result_col156[1] <= data_out_4_156;
   result_col156[2] <= result_col156[1];
   result_col156[3] <= result_col156[2];
   result_col156[4] <= result_col156[3];
   result_col156[5] <= result_col156[4];
   result_col156[6] <= result_col156[5];
   result_col156[7] <= result_col156[6];
   result_col156[8] <= result_col156[7];
   result_col156[9] <= result_col156[8];
   result_col156[10] <= result_col156[9];

   result_col157[1] <= data_out_4_157;
   result_col157[2] <= result_col157[1];
   result_col157[3] <= result_col157[2];
   result_col157[4] <= result_col157[3];
   result_col157[5] <= result_col157[4];
   result_col157[6] <= result_col157[5];
   result_col157[7] <= result_col157[6];
   result_col157[8] <= result_col157[7];
   result_col157[9] <= result_col157[8];

   result_col158[1] <= data_out_4_158;
   result_col158[2] <= result_col158[1];
   result_col158[3] <= result_col158[2];
   result_col158[4] <= result_col158[3];
   result_col158[5] <= result_col158[4];
   result_col158[6] <= result_col158[5];
   result_col158[7] <= result_col158[6];
   result_col158[8] <= result_col158[7];

   result_col159[1] <= data_out_4_159;
   result_col159[2] <= result_col159[1];
   result_col159[3] <= result_col159[2];
   result_col159[4] <= result_col159[3];
   result_col159[5] <= result_col159[4];
   result_col159[6] <= result_col159[5];
   result_col159[7] <= result_col159[6];

   result_col160[1] <= data_out_4_160;
   result_col160[2] <= result_col160[1];
   result_col160[3] <= result_col160[2];
   result_col160[4] <= result_col160[3];
   result_col160[5] <= result_col160[4];
   result_col160[6] <= result_col160[5];

   result_col161[1] <= data_out_4_161;
   result_col161[2] <= result_col161[1];
   result_col161[3] <= result_col161[2];
   result_col161[4] <= result_col161[3];
   result_col161[5] <= result_col161[4];

   result_col162[1] <= data_out_4_162;
   result_col162[2] <= result_col162[1];
   result_col162[3] <= result_col162[2];
   result_col162[4] <= result_col162[3];

   result_col163[1] <= data_out_4_163;
   result_col163[2] <= result_col163[1];
   result_col163[3] <= result_col163[2];

   result_col164[1] <= data_out_4_164;
   result_col164[2] <= result_col164[1];

   result_col165[1] <= data_out_4_165;
 end

 assign result = {result_col0[166], result_col1[165], result_col2[164], result_col3[163], result_col4[162], result_col5[161], result_col6[160], result_col7[159], result_col8[158], result_col9[157], result_col10[156], result_col11[155], result_col12[154], result_col13[153], result_col14[152], result_col15[151], result_col16[150], result_col17[149], result_col18[148], result_col19[147], result_col20[146], result_col21[145], result_col22[144], result_col23[143], result_col24[142], result_col25[141], result_col26[140], result_col27[139], result_col28[138], result_col29[137], result_col30[136], result_col31[135], result_col32[134], result_col33[133], result_col34[132], result_col35[131], result_col36[130], result_col37[129], result_col38[128], result_col39[127], result_col40[126], result_col41[125], result_col42[124], result_col43[123], result_col44[122], result_col45[121], result_col46[120], result_col47[119], result_col48[118], result_col49[117], result_col50[116], result_col51[115], result_col52[114], result_col53[113], result_col54[112], result_col55[111], result_col56[110], result_col57[109], result_col58[108], result_col59[107], result_col60[106], result_col61[105], result_col62[104], result_col63[103], result_col64[102], result_col65[101], result_col66[100], result_col67[99], result_col68[98], result_col69[97], result_col70[96], result_col71[95], result_col72[94], result_col73[93], result_col74[92], result_col75[91], result_col76[90], result_col77[89], result_col78[88], result_col79[87], result_col80[86], result_col81[85], result_col82[84], result_col83[83], result_col84[82], result_col85[81], result_col86[80], result_col87[79], result_col88[78], result_col89[77], result_col90[76], result_col91[75], result_col92[74], result_col93[73], result_col94[72], result_col95[71], result_col96[70], result_col97[69], result_col98[68], result_col99[67], result_col100[66], result_col101[65], result_col102[64], result_col103[63], result_col104[62], result_col105[61], result_col106[60], result_col107[59], result_col108[58], result_col109[57], result_col110[56], result_col111[55], result_col112[54], result_col113[53], result_col114[52], result_col115[51], result_col116[50], result_col117[49], result_col118[48], result_col119[47], result_col120[46], result_col121[45], result_col122[44], result_col123[43], result_col124[42], result_col125[41], result_col126[40], result_col127[39], result_col128[38], result_col129[37], result_col130[36], result_col131[35], result_col132[34], result_col133[33], result_col134[32], result_col135[31], result_col136[30], result_col137[29], result_col138[28], result_col139[27], result_col140[26], result_col141[25], result_col142[24], result_col143[23], result_col144[22], result_col145[21], result_col146[20], result_col147[19], result_col148[18], result_col149[17], result_col150[16], result_col151[15], result_col152[14], result_col153[13], result_col154[12], result_col155[11], result_col156[10], result_col157[9], result_col158[8], result_col159[7], result_col160[6], result_col161[5], result_col162[4], result_col163[3], result_col164[2], result_col165[1]};

endmodule

