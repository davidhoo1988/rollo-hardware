library verilog;
use verilog.vl_types.all;
entity test_rconst is
end test_rconst;
